--
--Written by GowinSynthesis
--Product Version "GowinSynthesis V1.9.8.03 Education"
--Fri Jul 22 14:57:55 2022

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.8.03_Education/IDE/ipcore/PSRAM_HS_2CH/data/PSRAM_TOP.v"
--file1 "\C:/Gowin/Gowin_V1.9.8.03_Education/IDE/ipcore/PSRAM_HS_2CH/data/psram_code.v"
`protect begin_protected
`protect version="2.1"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2021-10",key_method="rsa"
`protect key_block
H6EWvBgQuJF5yC8j2zjI/cBpMWq6x5YspBaCbXAKNSbm2i1pbpVIPOHhjfyusSdRZePEG1Vn0vX8
ZUA6yy4djKUKs2q0bfloMMjOUnxMvkfLa5MbipRC4j60kIUxER8AosLNt1ncL8J8CAe2BeBiWK8w
HD9UGBR0HgmKjneeHGgRbutt8/xUCfQ/lSJKo9aI6uJ1FjdMrs+g8i8lpuXs/He261KWTdcp0uzE
Gc4bXUkFa68p+FkwNTM/ZcBOSp/GohHZcXDO0k0JzrCRFsdN0m+I+Fzdy3WEG9TVygEGG5hXbJc4
nGVZ4oZfKpMI1uVyUAPC7S763m6qHbFs2foqpg==

`protect encoding=(enctype="base64", line_length=76, bytes=370480)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
J48fAtJmUoQ9lbLf90JaEwT2VxCUp/pf6wFq28vdpM48CibNJvNlrb41rN4y6mVU2IX1qmfMsZX8
oGJzb0YI2JV4IrYE9HWTQd4PYgjNyLwz6AozyS66kiKfaAWe3b7sfaSq8m16SbM/eacWUKPbyxQn
Faxc6jlGKTGiXH8BoVxA6smroyjaAgzVqzuPB/w3EJWQEBNW3OoaIAVz4L46Stke5vqfrO2qMcNG
fSBhteim96/G2+PFWExgzokbPUW2K2dn8bZe1digwm09BeyiB1GBhSNLTPDNHISjm5UaCVFAHO8X
UVj5amPF4r/vING3aoQTPgXwuFrClbMciQSCIpLQrNOEN6rHKL/zfihYqV1jL7pA/V0AQr6q1dTr
SI4KPZMJh3A1BWuVHNkeAJVLCGs8r0e+DJUou4QX/XdxO7YMzINCZJuS76GnapyoSKg1msbTg58u
ZgRycPggdK5Xpu7PbzaEfESzOYk4/6Ap9Ku0UFNgEbMtlJsxA5zGER66vyz8FQ2tQOFsLzqh5n1X
AqwYv3f5AKHl1SPFZ+mvgPPpg1EshrKHyoapSXuZBG8RvA1TUJm761MwCEMBoM18RBP0D+LyNXfr
no6ke2o6gTim4G6c8yXkSQPlJRXFeoYfvPBeSH5xhDh6RPgjHUv/cTkek4dust1MNhhQ87qu4h+/
Z6XloBDwAn+oYAxPpKiJkPRh7vVYSV3pYlSRE1T1cz9f8SJ2oPFyYWDx1t/tuWtaEiGV1V/Cralm
NB9LBE52OSfxB/h4uLV/3wEvFEELLPfi0ntie2OIJPLHZtuXYeexWPDS/drnA4Czv5dDL+Lyy+UN
mG1W+N3CAa3Ixyov35v1MzYLfVupz6d4qaRKWaUhqK3Q2/cm6X0Y4i2RWb1NPdWkR4wBcxQA8h5v
GlQi9+kN3Whl7+qfBMINCp45X/3dV9whPzef3sfQR8MsQBKDdjefH8cNtq0DJJPuuejFoabYdI9t
CVoyA0874Kce8Ym5AjTuzbkYuf9PkGwm4yQdM/ON2fPjLlsvsHz9KEnuiPB2ItzZvb9i+DGpUnO6
ySt6ZQjjdMA8lM6g625qVhCRQfW27Yv2oi8wjx8eYpMbcKCGLiWS/YfoCm3eH40ctt5/G1u8tW9e
uHGuh4UwyaP6+nOc7KBm1hZAy4qniNdtw2HZ3vRgQiUxxLCsPM4WnalGjYfTdzPZIE9NdTwAUtPl
hSdkQGSaTGVj8nZhlZ6Vl0KcYA5SJLcjzT16I3DnK17OrVrgn1APuXzlHE0qtk/s1glzaSTLAc+g
tLn12vVFFW3R2EVP1Ws2o2QT002qpM8qfvhmElcLq7oWh8FBFp416DECFJ+RhqraALpTrY1L/0zS
a2F/j8Bdyd8gdbreBmHTJSe32m+8M3Wx2ITQzcGio+4ntzD9hP1jPfDeptrmMiYumNvvSdqbV1di
IAzjXIJH7x5oCKcxuFC59QCpaQPYYE41b5dMGL94Ln8dBLgsMYvFDbs6AIosyYCR2zkiB0QBdDCb
UJuZjKj7evw+hJSrH6LvsKHT8EWXKDZ1p9q8SrV+3Ip4FADwtO2E5GFrGuvjOunYgVc+Zdtgt9gV
XEijW0p/cobwP2D3FlUVYEoFFidfAk4J5S0uEhQBYvWiDfvbzyQewbdJxjR/4vTFYlT3fO29H0uo
qQMTc4T1L2lUO0i61H+MNp4Tcaw19dyvZpWiDMlzrl52e5J0MR0bvO+gEqeRfZYL6tlT5PVNfzYo
1fD88XGe3w+PAxMfgO3Buu/kbCfo6bVyMmgoDx4TeHBI4WxYDqEy9qPZdxFKbsgYdQRsyHFkTbNB
JF2efQDUuh94RHkZEioYXnoTygiXURtMTPZzSWzM8OzaQfJDsl3F7LGIh+TRUzcn2etk5FQX1jBK
+5zfH30ykCzTnacFzIgmCCvcL/Gu3MwHxftYAUXsbKbodMIrEnFebRx80BFYEiUazbq+c77lr9IX
HeOaHrYDcDc7buOy2pcVLaQlx7663G6Y0kIDnKwbWMP1ETDi0DRYfLbzzGMubC+eBmTvw+vGcIGC
NNRmCtfWBTZaJVF/IcjblrryEM5b0tA2+Y2VOTWXC6QEXP8gXNvmGnSJyY/Oe2KPIHtCYYc18YBx
GNtCjyWza/l/Zg0eSI4Gi5tnJkl497iip9ABtnsrR/TpslIIWjzfZBI1u5VlARAjM045/sM+AiRn
89tETkjZfND3Q8ufNlzqeirS6vB3sbUcGyNvloQhwVWBEAaVXoUEcnhHCKwhsnNXNHnNyIwy2ZF6
lBXF4avzpUJyMzBHkXdT1lk85dUkO8FVe5tDU7qadvKjSgNxuluNALn1u1O0v4MwxgaCnIFepO65
FYiNNmUnMZZhFS9NmJ9dvX4mneK1NEdwZXiOGjzs/jfowIf/5hLxaN49Fi3ZjbOvF3fwW4XeTYAA
8Wvhn6m9VazvpCedKO6BdAFqbEHAVXFgfHQB0A53BRVG/gLNPm4fqqWI2fYnnisgt+axQv4VZNpy
FIKXAs/GvjdebHVzEhhJkCJc8sGk9nY9BaEwunI4ng+oQEs7rHcMLYyMFdnLm4Ugy7X28gZ6apgU
zXtGcGTYoX4N+22yvAr44SaOLfAnmV4DXNTGZV2YgIQ5kRRmJ2+QfWSZBeWpXQ8EKjUKg7KefQPS
lYqcDGFXePn28MAb+nNYfGySJbMwxFrvdMy31vOl73b2YdN2+yWFVPMdv7uTanYQ/V9ANEDOfyHI
icccaweOVc5Qm3oqYf7Sn9dmIQtLmvc25yPiO6lU0BeIIDARyyhq8hY1wrxqJ+XMBpdWZdEPPy4N
uH0Rxqe9qBatyqLRphS4GQsbZMVLr939YctT7Vwl6VY9X6AVHGQdQ0P/cK6PC4YNkGET4BQ6QTHG
br3Za79JzB+7ROPICi4jWBgicdNw+9ow8MkgryAVtXYco3m5rhp2+ri767mr7oioQWEmT+/Ungoc
7TAX/nC/EWax4Vy8HLemxZ7sPCVNcj9Pfg8JVBqLmgqQeJgmhiGsy52iJJ9D01KpeoorcsPfZifX
UYMk2RwwLkHBN5Xgp6r8KhgshS1hG8POK1nkUraW+ejtvqVY0d+ngrFTOX9IghbMrsC2aD1ezaTe
oDRZTKpIdwCGyRFN9n2ZVyyd5rkXt+0tpMQGrAO+hZ81UU1Q43RRyeSQE31Ycr0ldb+QpUySv38d
PLi1UQdEsHRFVXcirmLLh8fKw/4FPL43XZ9DnnJt2C2wIp48om+8yytgubkSIooPhgENdRZrBPLb
mDZbjcsi3K7nU/esghdybTO88IFccHz9K4G1BIIhRRD73U2fKxisfYZEihD66rOcXfnH27TPpwW7
0faDC5PJDnAch/WzK8ZUE4di6NcHji/z5QJGYJFGVq4p7o9WnrIf4198h5yS+sCC1rrQ3jm4nP0m
0W4kyIcX1CPhJk+GfZvbM51ZRBA8bEJhiCdhdlOMfsfqd877dxHMc07aiLL9WyNvLlOUaNxDIQjG
Gg2XVkBbhEsP4N+Tq16GuTzyJWWJ3i67MwBnnhRJYpIiYFsUCCKRPlLwtmPqz9odehsBLCxzcvrC
LJ49IVGWFK+b7LudNFlPAKFKw9y+ncX29ayiJbN/YDAVmioOCvKq0D/YOrFXTuVrKQfi7af8Vtof
GfI7mJB5U0u9Tapt0oTrBY1MrdvOjGzFAy7YmzHHgT8JMXIlaMn1+f7WKj0Yb9LGTxykSxZuMY2Y
p7tLqMdRe91AQNW6bA+Gv+i08WHCL5evJrTZzAruqymPeaKkh4RvNG95uHPB2AKmthQ2uoUMaai/
0UgJedZdjjSNhQqXrHCaELtSMEjT32stT9r5wZLRjtuUzXl2JPPPqFTxvq01aCB1Urp6GlkZbkgg
iSJYAv5M958h6ZD40W4rfUid4U1BK5/VXqLlFGUlPCr7ikLT7rzAod5YDD66+5Ze8YuWuAUE6WBD
mkLsti0/K7kwucGPZQWUBAZS7UFvGS5u20hc4ASLE5lRc9d2y5x2NgU1rBOQnpZtbPVr/BJOgiFo
lyE9Ra9Ui5GErK9e4yqBgnGiyHUU6NwCyk4GEXIV2dwQRrablykAUdybwImxM5ZIXc1+lx39ta0a
bxvmrlM9UKLVTLP2wNX0UPBTfx/YpiZZ6B7CKMFc/daFPUXJ8SL9kpXlZr4jm/E1fu8hP/CzdyqF
juzAXW6fqQoZZrL0LxcoOptWD6gUny4NySf2F9aY4N1KeklUAj2tO1yAbd70BrDoCmrxJwu9B1kc
HDKvz0Fj7CLJQYQDb1iXVAmTO3IOKYFwBCX+kucUMTNQayaEgx1SPZdg9AoFIEpm6JYGfhO9D8Kf
Yed8GryAUiX2uRwvr7+LloKfoEptUfqz7MBCiuFOfQ5z5HbK++KJsMi1vLv8OYqv29LgT/j99OxW
RmlaPqVNFrRo8wXx62SO9ekaLkuOLwWZZOWyzwnMEZgs7cgUrzX7WEzyD2/XwlAAGS424sEnbxJS
I6X/iT10IznMitfi6ZBjSJhC70RA35E83xroD/nTdpJUSf9y7QjFe04tMr927y6/qqlIIRl+bXI8
PU268iVb8s8/2StDJkIYV6YyS65e4ry0lVOvhq4aV6dPnPPxtE+lFEMLGVI8YTkIdx/kv3a5E8W9
Joz4VqS0/cJQbxfBG1B+ZbveoZWTJFmsvKJ93m4jBGJFuLDx0lCn1D8VOCtU4bvKTiNAMxzO55ei
jf9378k6uhQ5Lht+xPVytFiVLTlBrYp3Waf4gMqqilZhZO157+44sZoju6/nkM16KfbFlJSSFetC
1rNS+xpBp8h2qQq3FN/OKyA5jtqjL/k3IzPieszolAn5jIJqT7y5hAS5gJH2EnEnwg6ogvmanIZ7
nJJuEdhLiKP+QPLuaUCGwWWQkpwzdRI5wJxbLosesa1Ps0ngyf7gEYHu/EviDsLYzomJbg78Tq74
qt7GkcHIhc28QQKupr3Lr/lLlHmoypZIStZe2JPmCtdf3jojQE04slx3dQndNwOLxK9VIwanEQlZ
gq9LyDHlq2/0YNfX28Ow3MqphcgHHqowKJke1fc6rnh5DzDyiKWZrTrCphuQwHAXFnVFiXWydKeD
tOZiznc/aHFgjoCgw1VsLIP40+gw6eqzBetB2Egux0s8alyXa/EMqlVefKRjFAXKVMepUrsljQUz
3hPVcMsH+T/Q/2z+iCBOmHV+Nrg6hjxq/+ccWSdNujjvEHdR4M0EWtznXHKLoRpN6y7BodbIS/7q
+9J0DmLfZ1dPTMtLFV6ES90qr4Zj5/uh3s0FgXDLBs/rljuFlXE5qo3T1IZSL4hsYhj+xiV4UvDl
eI4et6vo8zfUmuJenGBHTiGxUTH7Fsdh/7XBG3oSqi0gTpMk6W/m3VeFAgNnCnBZ4xey8SUn8wrO
UCJHYd1dhRHvht8mLO8FNplZemJerwE+xpYNQEacsFKzZ8LSj6olDW4JG4NPW5vxGgVQPMpjm3a7
CLpSm6ElPiguFISOL21B4jDF2OhoDsgCZ9WBDSfHE7pIPS85CogtNIL9VYmj7aK05a9Q/lAcXDmG
PVFvKd0wUnOO23gogyirC1l8ZcUhUKqKM3okp2SxCdDqPiOqxG2sDqBfVZYHo7+cOFnc69yAtnYv
2PeXCtMN3XSnB/sdqcdvjqrKhZ/79vTmABnMO4tIZGaA+gK5HA1eK8yFaTwBnd/IseMRM42R7Ue1
PfYbqcXCqBC1zzR3/pvBjH89AZZpV7tlXLtLHhU2q2s3Px2kvXl6K6P5E+LzlD/aqJ/MElcNdSY1
nUf656d6wTsC5QGzr6sLHRbB8g3PsBUbbwcWjlRWIhX82N2UkwR5fi1KTaMsT6C6o62wnaEyLFpn
tE+RO6ieQ3fQ04HjqFVg4A+52UXfCTwExFvzn98uh4FuWVBZJYVaDTNMEdHWjkPkEQIb1RrRFAm8
TbXOoMGbI0l+rUUEFgH6obqmOiNIRPIsbo0u5lFtfW0eY+SDTAppv3cYfHjXeOcNvPtCLxiQrFzi
Dbrtpd+Rz8aFmO4EVpRV9wODQLBK238b4hT8YjtCZirSWQ1mb3KFspfncRCeoZQUx/hAKAvwGSNl
BF9O7dswddmgUhI7q9/Z5pOoiKh+59HRdg9dnSJGd4t50EMzq4GY6KpG1WLHUlb1AqPUbv+U8K9V
sDW73T+I2mm9mVmvMIRkBtHOhvTb/aBBF2hwS5DLKeUbX43xxrDZSRLAp2tPFHl+3sJczPjENQlK
nx6YnCagWBMZZGKPx3HNU2a+TEVHn6LajpsiCLpURTzft4gax/6ax6Ds0y4nlNubogsRSNg6SOhS
V2mSOOx2N+FjcPah56TPLgm2Ssycmcb0C+X58BzGQd58DhgDV89E5qV4nq4J87IjRXTrHSifzkjx
a+9GWmgKNptVt/BozAHwDW7tLPxM+RSa0enTIUM1oqXC+8YMoIbL5rTVFHhEYH49eXqU/c5Gpswf
GqmlRK1FiGsIXDyRcREWrNPE90owLxjkmV9jrtYbYXsRjNplUeWKNX8GbAmjNTLlDSyzhfxGlxMX
wo2SCkPMrkkQrPPXdgVAgKcbibJ5S4ASP2sbha9rBIQNGhoTwzdXRutpuNlNyOxquVNbIrdAuBM6
RhpvLEUD4Upg7Lo1zaCU4uajDfkzcfYyDOHCeJ4vknS5/HS/T7/Lu8SFQUNeMIbdVr4KPociBiQ3
pUnROuC6PXtmXpMBfw3FE6S9drh4YCH3HvmEX6szw5+g6PoRGeeCS07q656MLTk9lqpOea+SxU8J
PhsowSU8nZudC3P05JvkP69a+7U3zhePAwZO6ZFwpG8lIJs3ORJEJBPi7dsFQo7i1h/gph7XaR/1
Vd1BbJT5Tdz/+xKF71pwBvW1ZJ1uc/C/8ErV/4I8XnBadaSfVci+ZgLda59/zNiJzDR/Z60cbTRA
4tlIYokuVup+Va0evZ5FwM6T30bntvf+Yc9BF5T33Q8tOm/TRUO3uWBpjeiwpBlf1aXT6letQB2m
q1f1voFHSQQAIeRok2Cm7++azklh5kUTd6BEXjn3gzXgHL8mtiwYnyC5ZEonPRWiA86tWsSFRqFK
wPxO7KCVpboDcBWMKp8fH0pXEnjwQnXIt/WJzO/VcEAPbqoLpBGGpjRG10BmjrYlAUf2tVZqGiTI
wjdOau/IOhiiPPFMQoi/xGvPmTcGokv6qxe15RQW0vY5TQvOnAJA5u1LcJWDTzuAo86iugPnU7f1
dlGR1yaeffBQRYQuPiRGAzftq2bagBrXa9th6eyYaVE+9MkS4jvw+wmAeKBnATf7qE+nKQfT0kiR
93JGPs0uTwzQnnF+UzNu8SmTyjUwLEn5vUH00DjHATGlNEMnH666dQF34W1+M47hiEVdsaVY8gMz
Es1vTNLoGBpLIH956qKyJD40p6wpRg3iBdFBSyy/Y2k9tGyBChR+QSFJXp0NeRrX1EF9Z431JTAP
vzyBksux3O95f7gbIcV2HbwdPQNWCnctmaBFARYKwjSvq/IsiImVJx4kF5SrxN5keXROIb7m2Kmf
JB5izmRZCLU552L19PgjYYAadRGeNJmJ+9Lrj7AI65NFxo49slw4LNtUV1YIoSBLzCBIw63EckVp
+LTQS6nFSD3O7ZAodg+R2u9pT7A3g/QguICZOmNuoRR4sPo2zQMLhD3pC969qkWsTicuLLU+ITGY
+Oh1RXV8Sp8iB574qqIQ7I2T9cGev7VBSZmdzSf51Q3tnFo/RbjBE/ukj6o94nV3wmNdXdJLhqvb
9SzDNjBHBT5USo0vj1U3bkJMdF0ruACLV4fLt5UxjJykw7VNke5+TRRLe7d5PgsLXGj2MkXiZqxD
mQcVKH6Inj9ftLHhJ05YYR8tx1r1hVxMtBEGzEIFQC4j0hxLjlW0CMRFpjS3/L8IYzkVXSHPwXRZ
aEpy7ttLWQLmKAOxUMRE9FEnFEeJ9Ejd91DTp4r/O9rmvesuiio2YDC9DqyDPtxFIX+XeRm68S8O
tyhK2dwDTNDSIlCnjQ1IZlOx9t0T3WU/ZWm1y5psHDc5Qb236Yyo6qED6aR/tIipBbE4Tk0fEpwj
wezQjfUXy/EAoAuA8ClXDbNBJgYEgHwN8w9gOGgq+SeqnLyGopZaAAMyV15OrcOl2Nqq8wmohFtb
7YVkoQ5Hh6EUhQEPBpSfZ3V7Mw6axMxP8HZWGbFnsOU0xTy0X8tW68TKB+hUHhX1AQE5588pU7lQ
aRu2YzQiwe0FJ02iwyzQWwdpm1O5TRHZbdyv3BYQ1LR1d2m5B2uLyS9ybRotTrjQPSLwpPpU91kG
B+rv5ANDdra726kbr4CZr0jOAcpufapB7p74T5vTk4ZNATFtip9nDdOiyQIyR6++f/16+jHnAVlM
KFvy+sCy+JNQ9axlO6FhkFvrl3JT5Y7tB4h+zLr1SX7XTWtPIbl/l0hV3A7vZyVjvFsfM0nwa1KU
/gjPSZyrTLSdvPIxFQMEwRKYPZ+et9NrLO32qKA62nrSqeiMu/AsLuEqEN7i0R/9T13aEF0UlwUa
kQEMgPpY+mrp8LSKp6tpKFkXavAYf3o0ePBVrSKP3FVW+AefWM0VIItlBhxQVZW33Hw+Jxug/t/g
USxS6Kz7R/aBzutX0bLTfxg2sT7erR1BOCHB8A0PPPpsn6F16hiN+yebkXDGFF9xA52qceLlCzO9
AUeqRwh9E4+R2PTqfvZCHx675CZDWt45DV94xPB0HQoskQrcx9BBoBwmJNhfPx1Xce0aHybMBLBs
oVTJAuCysnCFfp/bbTVPQcRVbaMZxX+UZBV3KmxWHHbVItNy6gu9chUIdv8p4p1muC5QvXbJ2Nm7
stc/wX1DxiFn0zl5f0ZEwlQg3+4e3faJtIPn5U2Y4T4iYmOrPyZ+cRPU9clctPCnVUR4ldjNiZbW
wIqbLHYeeSlYw/aZLeSPnpe74adExSfO1OczNsxwtk/S5ehWs7fNrqvz9fl/xqWhbLOYkzdlhTGi
2C3VBGvO+2xe1+6BiW/o2L8gFrmFjSwxWK5aQwEaU7gkdjko3GequZZfN0mZ4Z8siiw+qzlQNfnl
o7dni3Rzk1GeNXGbl+18Yek+vdJpe1BuYXjbhU7bHn8dxVpVr6oqXv+TVyiM2Ha0cIzNoPnhyNSp
gUZDnYu6q0ycVqhZ+1v4LM7+FC1XwS1/dbiMkbyuvu7q9tp1BdUKdpDUEIktrFwYZTjk6FvT6PQK
1iF9YHiEQz9kFtkR3TiwFsiH/OPZ6Khq/rokHcTV/0nW/6oZI6rCB1rkFzBU4kxO4zuuLfqMU81I
fKZgSmuaAZtGhgKkn9E0cX7XYvxLOIH86mrxqxfmHaSredpH3y7C1tKwKzCYGWh4ZjWTBUwu7HLy
0nej5JBSX6pdmgzNAQZbv69lcEfD/eSScbW0XYqze519g5h9kIKGjqSW8hDE2aIElzstBJnazSO2
ANg3RyWrMmCE6J2uVTZdos8N2L5kElMw/UDWHrYK0CikXoE7u4Y+T2et7+YrIj2zVkp4waHMSAwY
t7WgjyB6BZdkxG+r09TpyB8js8SRDShZ5HPg6qFq2lF6FpeVKYJaEGWCXQI7o5dKn8/fm/hHCITD
WYNgD2uvCDwqEtGU7WqNuUOLqVeT+dKRVh6vkEHzwO/dAsrvv9Og3cCeHI53uIsXSZx42EuQgTOI
PSftqkIxu4dR8AGLkdELTOz7dwR3IvvqdL4IqBpCDL1vEkI67jBBIRGIHpMFv7djhrhbqxCfAhxP
EJVP1Q8k19/CztDzyLYm3bVId/VSwFGR79vpsQCZ999BgivBo6JYTuTtO1HYrtcYlwkUCDAIavcw
OMe+yDgHjIXJdzWgQzpk27frV56dAWggJFVvw5fwWaGIS2Dx1f5YFeC1rwCFepdj1CveK99E/IOK
CtGtVhnxw0rglAwpNpyvB3dlwdDQeWhJV1S6jRpE49WpZyYpcwrhHxH75DW/yB/9r9CDWs2eXNqc
ZaxmOww8DPXh8ViWZ498pLmq4sE9DPgEjoo/bnRXRdJ24dO0u/NYPyXpPat3F5Oncs6awsWB9oUB
xdybMmh4NpguJxzD1W5+ROJ7oFm8KThdh6IH2wS+0sOBt0QHe1ZdhvXg1NTADdTTBD2zlYiSBxMW
u6CltAvTnH71Y5g8EmFhCqT/cabVwX5dIUucAo0GaHwMNHS9Sv5aScuS4WOvQvjHGM0KAKim9Y+p
t59b3i2r1fZ093nr4AMSX+EQpGIcO2qfiAIeFs/2m9Z5pCTcyvb+W724Ssf4AzujQt/g6yvRVgVm
X+wGaRdYvWByw9D6eKCmyB9mdTrRmovIvsTXJEglsJEp84EeDAgtpPRxYFlZ9DHy5TDKLOo6xKtF
Xr5hAU6o84b4sEKZeNk09WPecYc5uFldJ9K1On/ayws7SklGq5z4TEGMnc9zVBZUfSWwfgqMnzB1
/LvZIDmpZghiVXkS2oTiQew2c/GvrlDWl77WtPvni+ymC0z0guLH6ZhGultEwGxuc41SSx0uRkHa
D+8BH2XELf5ra/5V3KlsU36yawITSwQUvOhylwgzw4GCqcXMaHosUeFrKpkk7jlGfzOrmVPH6UY5
NfP/EPFeZVqn6z+FHWQVXeBYfFrueITxxmndvwDlHnZat1eUukJVu9BtUifWRrd8249xUIBW2U8e
mKYYOeHHJTkbe4MeH37qi6ZEnD/TA5IaYJ28jqjK5QnoJuTgWrYxeBbDh0rCISg6l/+pRhsyuU6Z
vt9TRhLlQvcH8ttIgovBBbcw48JdB+oPWChso1Opo3vCE0a1N6eTNeVD+Aj9sR0w7/bU065Dwfbo
O00v9YITKY/BZJW5bEAWJ6Ljf9SUD+avE/kuP29xq90rr35iZzKrMFKqy7/b11L1VbeyRVO+t9ib
+4vCKD2IR/QxYr5aAEub8Z7ZxIcUTqPhTRAfHg37WFp+qu0MSGl7dxQx1EdSDWq/AAl2eJfnQuJB
gKwZkV9jHe2e+rN7aCGE9YzwUytRjPmS4iAr9KTJenoW9YIHLEMLpqXl8PjgMlIJi65uvBJyeluN
foavi6NQoHrcc5AhCLxYBXB6h5DUooA4r1g/SsPHPWjZV2Q9H0gXxb7NZ4Edpd3MVvHt/z5dVwwm
E0UQKYW8t/lZzChuIfPw7juPQ1qoJq6zhQxRSoGcAzK6nYZlynvxQGvizlG6O+j6GQzdIm/WxWz7
IyPCf5c1Qv59cr/1NBXieeCUONnq0RmoMJqzeV1zIGBoESCEBl9gGKdqqlXtk7zHBupminbg+uTR
62YZKbzam7NuFr19s7oeaO5bkItq9iObIgg1FR8PWfoYrwVQEJMYxeORDou3s4nR0vFSB8NQMjCA
5id7Aq2FMo7+DCLBEMqvYCVLbpoPUvdXHUlsoXRmpp+PK0RAkEvqgWFX6HjLF20RZHTYr8qPk+GE
S0KJeGIdu8YOLFTj6pJxqeKHpPBvGLlMd550PmvAtX1sihWOZGoa8TSY2A7s/CQbMQdDILKwtGWG
/V6k6U6lAHJgZ1dZ+DpqHCjejf9CCd6mf2Xl5RDQZlkFqPxtOG9HShjy05FXrNH7fj4H82K1lCcz
ebA2Je/NITWT88/kA7sHF06nNzxOVeFVfXjE6pZNBZUZ4Av2bNJiFeB9A96QISnibj2FmaBRS7Ev
q2pa3E/7iWQouI0oZWxY9egFjaJ13RlxZtQnUO8WPjNutO6TMvqOkLvyvhCSfX5zX5JXqiTnBMPC
sRWHYoarHXPaAcLS/S+tZHgvcKv+ppaX3nngieXP2wxn0xlrkxSO+j2w18qK3QeaqcbIfkW3JcF3
0iUGTh4Leh9oUJ4w1Gl8Bgk2u0wmJgSkMGL9mzof8v6QXCz0jgFrjfAaGpC0IuUmNTrX5VbzEvw4
1l19X0uO12qzKWR29fvzRD7Rjw3N7eFrOKDxyMqBNor/duIj6deW88a64eirRXwUGcSbDSaG7aJJ
jj/GW91agk7StkGPk1+CGp10mAJqPe65aX6d8FwnoA9wZeIWVsR2xJPNWziZSPEIWX0Ev5+tomg5
VCD09ZUq7b55995nRY565DdfIiNg4bnHIFKbczAWT9JKvIEFsXaxKOKNlVxgF2vwMLAARACZXP5M
F1YTmOwXQOD03V7KH7mzvoWMKnyKFJnyYs6RADxj998ErSfXl/MCuaqxY+/Jk4b4C+IC6gJBRzAU
zerFNpAESXBTVc65ZESndsOt+SoH/N3YPYaIkKI1i+wTbKjisfSSUjra5f8hwFtR1wajjt5dkrgs
y3BNUe7RRAjSEdMmjgI0ycUxMRGjNIsu7d0MpfeYWCRpAx6KjivsnUkYoAhm+zOuHjzD6TD0kC5Q
gP0Ird4UuTYHYN0eZ19U3reN1Gly+ZN24rx8ZvZ+uJv9cthUzYfeopisRjWxF60q8dcm6DWZx/Dv
nOvv4TqPISF4SgQIKmotZISygcrCfdSP2f0FK2hvkvNvF0tsGwT3K/BrR5J8aVVyAZPt2o3tvAsC
Rh0jljVyM1dyHaXnYP4OZphVUYWwdup0dgBHRUPwLnKXXsUrhfXS/FToL+VLWpX65XWl8/nC8VHr
59tPDHw8VDGON8up85fvwAbQbnuyXMbvrWtxiaACAzMNMt7cf9albuGKfaxCoQPWloM8lXRm2JfD
2EppwqaCIjKFUwB6aKl6ZZWFB6XbeCLBmGXER1wg7VzbkMoI2rR75dSbLs1oYbEaKSdJUIQgJdHJ
rVmCx2mIwKKeiUxlioK3hODopDXRR4S2/0J8oiFoYvo/YtLiry+7njVqvR8pCeK08gfvA07ElhCc
DCPL1AQ8s5ft3GaymyLYPNbM+KDudyS7Klr3BG8qomdg2+Mvo/c/SX2AQt71dUAFZlk6dyesKCFP
QeWUu5MigGJhUr0Yn1j0YTH7hKpiapGblude5hw6C8tLhIjarlMjKoA7Bl+cJPhdXOZoIZ4EgrNP
CSNa60Y6F76tuP5oZUY0ISz4vTTbxwD7YU/xD254wnOEBHsHFCRVJxJbFrVVH/qF4iAwEKRbakm4
Sxd3cFHSv7jLmZqtK41TiBjwFBfATo/jRh31mVwJXhgE7NNhNXwxHxmCkCOT1azmxfu8XLTL3fXF
0IarOiSLRm0JifJO4mKD5Fa5FBmZ63JOY06U4j3vgcqBac2jchgvzBivw3gRVZeEL+e2nnIOoH48
l37AY2fBIDUMJb6P4nmBByBNsSRpSEwWMBImxriuJ4sz0TvPHFjGUBMvqW+Opk8XHn+Vm7Oxp85R
BYr4EfAeL4r0NbWFlQrdsxnM2qY+8JL7Bp4bAqcuI3lYhANVX3xwmbmJxHenzK8xIOuDRHqPQwrP
HbzkD2SB/ImZCRYQpbATAMouzmIdF2ldHouoY4wUPbD57eN5Wk8ksXxNJXUSl9ySww74DHkn9hSW
186Yi5fVPi4zr3pONS/DnJ1EMrnMp5UsrrLiaQGjpv4xothVJcEbBSPIpjt00QzIziqv6dzaI0Ut
filyE2+23dJY0J/k/c1bk6eFQDpPQW0WGX7H1ii/6Fh94DTBDl7R33F1tcNncWLr/hNQrKUxT13c
o6SCHAsMSbjLNV6c67/XnaXUSctZeWoAyDBPiSgR2HSwPEJKMbLjS3J3Y7LT0QJUUPy7rf+htjb7
JfrSw3CfZGmoK2lb3GmeAg66BquiGl0bD4rNrisZDnqiIrdGEr2wuT09td2ekkYF+qdSkHunn/YE
627PWWB1dAEe2xwVy2xee6DzEGfKsXH48p21jOjCB+n8qSsdfHmdfNf2mW6rBRsKDUZjHKBvcZ0y
h4dq3/xUPtsktIoHh5I85q1qGt7FYb8DHtI+KsasQUPZnKsOHphqFMTe9pgPk+g/zx5dSmVymni0
P6OYFqWJDe0gTXr9jAtvKMEVxPdkBriYe29OtgLrLAI1rd0hQECqNIBQNFmSOjFkE8GVSirBA7hT
wM8yOxKBGyXuoduaqyI+47UAGt5cMWG4L4dSD911B/MVsr/mkOachHGp33i0F4sD9JbHO1GtkFSF
brlnyAI4d/I9UrVE5hfRCmq4eNAgn8hXwfSjEWDI2rhEmuhR3gM30kfCh/gFS2FFb2v2JRZgBrGR
Ivn2deSz3sCcCaM3f9z4YBZipHv/Ywa+ZB/HO+DvlkoaCvxZWKhwvUjsmBEYDv9N50nPls+SKyas
MsJteSCMC2YKO/PX6Bw/GMKOV00maLFH7Tb1EHCX5YxiHZn3o+wpMWrhDyf1ibnTBweTRekEn/Fs
Lmf9HMYuwEbK5lNB4jUHOgNWfNIwgeoByGOC92jZ0787HXK71y2iYDelfQatb8QIb0YoZCT8k07V
COwodFwZubKjqLKM9xhvH3Vz1fNacVO02XLthBjpqjMB5kmlLlCWlW6zeQglYUgSCjTti/0WHINy
7H7PFH955R9/+dXZIJwtYUieaDPhok5rqy2sL0x5A12nJF2VmXO47viY+ICNU4EHhv1DjdXmu4Kh
wcS8pLfQf1s/UWcezcCYid7NOS0aDUYxxT24co7z7xbk5TXcj4IVx5wxjMnUdLdd6tOH/gDDCGE2
Ls5mS2FF2LwvmEWIg4lYbpTW3qMbNOslV+dxeY2HDcsO9ULjvH2IO/216lW0BZ9m87Dmd1L7N9eO
M0mOo2raGVHozaY+ZcHpVN3ijrWfNN7sUX8yTZ56zp/RuUO1cfntknFiVWV5hCU8PN/bGgD7ae9R
63mt1EkBA8yJ5Yr6jUvx/wfnk/reSqb5wIxhu4n9OwJAEuKN7oXi9HP7sXkft1dbbXu1xNJkV5sW
I8KImoalT/CktoIHXSwg40R+nzZzE2Ih4gxQtMBTMZ69YxXqrpqKBBFormEbnj+I1jTHIOi9veGQ
Up15N4kVK7fLNwYQLeDIraBsLn+BQj3CDcHRLjwsaWvfmHmMTIs34iijuY8pdt/Hhwn+P31opUa8
zdKXSvq+9jozGM7Z5Ly+YkAJBDm5mDZka8qQ41tNrbi+G0mU/Yn0m9DZkHsL2J3vf7ulrMIL778V
zNzwIXXGms9sLcHR+I45aTeYUHkaITmiEqVe4cnky3u9Cvd6h/qKr9+DjJyaEFJEFVNo4GuuRZ5C
fFVxdGZcKg9ziq8rJi5sTUfk0jtLOCQwIzlAR/+eYaILzw65fw/O2xXAgEPpS1YKupYpJmQ84oBW
7rI261MvjgPXQBtS1rzDn7QEdjMH7UztzvrJTFVXFDenN3spxSHvUpc2q5CZG4kZ44X1QzxDIcG3
hgZRfKZ9eyyHptYNmpoxcaoTfAzNG+zkjzJk8I1gHqIcfEqvKVDsOd1N/a95COArQAQYwR2MTMrf
FIlh4fFylPyUBCuVYIbqGAW9SXJVknTqDUaqOo/2i5+adP+b7xDN4Z9kU0iXOP+BLDYEYrxo724R
yuyr5MKjJXEpbJmnH0VpJuY2/1EqjSuCfTydAY4tgy7wxU0OmP2TT0Q8+teSDJ62CJ3ywSdWOXot
TRAhqt+R+bjL3hIxHDYhimV2hagxdj4bh/WkpBsYIve7zltiQWX+QNsw5Wf95nzYVgDYPQkLTNha
pVCXHlqS+NtlNMG64r3XtzpL1d3m61TRIN5ZdHPcBeByt1JF0WqYzDCJZoy6CDqe+lSc1wgSyekq
ejhiWUesK1Lpn5JS62Q7/9GRY3LPyU+v14eszs7dnqkvxvmCxO9Le64EdqI02wokQfYbMqVIz+4U
WMaGniLAKgPYc0HdykUK6k9bYhkQBucUEAWZvIAfSDRA60SAfsZli0+fYivSAuwQponF37VkG2Df
bvZUiCFnuuXIzLxHJwmgNWam2V55CI2X9wMNnP4kPfy2d4hX/v6gVV4/weBHj++/6rKke0RDmkdv
PCij+jPw5FJuGtxUjgGUW4/geKCkBn+qftsphpcDyu31BdLx9/De9AVxEOImbaJsnMtU3D/IX4jW
dHNGPRNQSAn6v9rIsk2XcQPekkZuKL5m/mOr8wKTbPgB43WkaZ2Bg7abrkuNBO3YTEYa8P2gWequ
ysub0KDzzxclItV0zHKBPmTrHZO7rwsGi+yRZcxkofr/EPmjuRTw2kze3/TdOz0FwfFTHRsYnKLb
OX6XbXsws6J4e4TPd5YZuYQ3WgOAWhfxkglFQzGCVBn6+PIwqWO8yakm9wkUaeknwfXhTEz25BaS
9bKdNhvUAPBYWfWXUIq6V59TvpoacGuhMbEWxL/Q3V4M1HSuvJOAw4+y1JycAvrVwhVqtcBbB0cU
u1moOHGa9wiMsB1MwAjcyEL0nfBi6NTQtohubUrhFDFA4fwmygInXFiborpOTHePxSRU8Rz2pBjX
XkwJ8t1gIcsO60bq0iaaVoERcW5vBnyVcvIlEvfAaJ3LCXoViCmH/OfWL91xhbXzw83yV/b52fn6
4FnC5VwZl/7ALFMEiD8Hk/JJbZtN5q8BYPc24mDspiizsV46W4kfUJKVJCegfPybP4GHYUHctd48
zM2oeC6fDSrhT5k/2skrSNWw8UkfSs2G/lnr1NTzzJ2KNP76SeA/+v6KWhiU84TW/KDguYQTzcaR
3aL75ZsgpyTslWRXq1zP+E6JiAWFi06B8VMHdsN5arvs30EQN/eVDO8wSKaO1/Q5osTz4A7cj4U4
dSu8T2Oh5Cq1NVL8vjoZoZt8hpcHZiPYeS1aBZO12Byzs3lRZMi3sG2IYMuCxrXsrrwgeZBpm5bW
L0+s+kITi+LS0UWksgrjUJ5eJ796pcevthdJkZlKmx8yqYlwTZdaElmQyIQv5u/Y2REJSZk42l6G
u6n2NOkgJl2eWvkbLm/fNoASpC6yvORKEZQjak7sMtTdlpQF7LNE8UwALlz3QtQ8sEPpEvE7ft77
h12wUfz5WZyEYA+FjirAdf7Ng8U1iKHfSvlXYOyuB6sI9UYqK9n57trygE8AAQzgDlFeoKuG7h3D
m6pCZ8LtDFqhsYYyJw7law9OLzUt7wqgfsoytNLj6Fmdq7cVbl4Nqvjce1aUqF1RWIrAUbtPvzRG
ZYzfks3VUz5ou9NX092fmxkbhZD0APQHvdj88z82/6JbHJNR/HKDJF0fpB6RizWYFWAIgeSdqFbF
BbjTWMA41p0i0jlFHms89xP3uFL65ESpg74D5kwGsqPUyBxH24A/b59kqHsbsbB8g1JtX0ZItdHQ
CkY7yMVwRW0rbx0vWe64lWgy3mrsKdNGen8R2iitzOrFu33W6j1J/hE3xMZw0mOSeQwV5cabVC2k
Y1ltrBOVL9vpnQSAA2jwNGBCsSrJNXvIzdQJ0O/1PWdz/zqPVVMte/TX6gA6mBE+t9SLroHt+ZX6
e60dHshtV053SgoanFCJqqTbyvIR+ukbUAKSDoNZ8Q4XvB2W3UjsO1h7L8doRa3v3wKNSrnv8n4u
M9HrjMHnmhX7+D9i3AMqkzg2+1Mxnh8MiV3DqjP4PkO1qUdDezcNZmMmELoU2eMgdI2QunbMlQDL
r1uzmgyrW5oK2HrIJXfMMgTPi+Y26YO7aL5bwA577pV9d8otS19fHkK9c7tbn1ZlZeZ/QnbDGh5v
4lcWcjTz1wkjmNU+k2uR9Y6qH14ztKmVWZfWhPkjykXHrWP1AcsbXBRd11yvdl89w2BD/Po2TYyq
b9aR/0rI0o91lqO236tqBhTNvAHo1nJ8TpHXQtLxbYRdFxSzRJ8BTAlzXuMPZmimttWiiC+IhjWU
v42Fj2hlp7qC22YHSzXQsYksYKj6fhjJm42WQsUPKdO649RJLsdUaamf8l1JWUjUFHty5cFr5yXY
UAdGIAllGPLMAYltyXd4uPNlE4neB3zVaJep6RwV91qVj0WzZL63Lf7udJI9b1UPQ0NsZNsffahE
qvZ/DpYVQxlimNfm7ne4o4MZJ7tP62Xu2J1w49NRxwyisqUDcCUOVFev4gg3U5qvp0KzUaOt+rPx
qdZqZ+5l+Us4fVMZnuhDk694bGGlWdNYhLBDv7uVF/EB4tR5OKK/pjb6U9KiA77MG/klMvHn4EMG
LamuxbebQHdAym/gN+QsqF8F9bl4BDmKqfnnR5DXlhlVONqLjFgLHGu37/MNp65wYc8ajBu+5oV3
VX184h4ziTKSXMv/eLFOppzPRHy44XMN8lAP/Gyzbp5JD+YLQcIEPDlu6HSR+8FsSJ9myJRdVa8p
l6CMGIE6TpjlfMT3RVQrn5ZGsbWJw3aIY8Mgs/1OhsaFniH3Il4kVOpX0lsZOz+8cXE72e9KEvy9
8ZTrlYMLkYJL+AYv05ZH3gRBr01KKn7qw5iMXlkOqX7cnBUdZNPVi7vPwGbVV9pUBbdBway8sfNV
E7Ni5qJ1hvsdCwwqrPllIfaGtTHFOo5UfIuqA8GR50CiXR7rD6TozsCGkbYUfV6DvBZlMz2/juSL
1fJ+HsGk0guxDHRQcvH/02PC64mFmwsMeVWiVkTdV9+8EKr4pUJOr/2arwbtB+gRljN3G5JSktOy
1k+diYgAOa1PtLUkwWbGTfDtM4V+cvFtB7hI6P6FBW+wL/l0bab/zJDCqFtx8POZH5OlyLNoWUYw
3jUkk+qZ9y58Z8kiNkskGY9AIi2hg0tvOE3SaPzdbZwXaFX8BFrRGBa+HK7AfyakiA7oTFCz8ygc
+j2yb3B5ydLfNR1TNrvy3aG14G27ZRhOoriCDqcGQECNeFSu1POidQXfZmOBkOhkEVRwrHX4GS6p
mXsjSlXVdQzgisOVIgwwIjaYyrqRfxrHtuLxZn21tsnJsUyp4GgBeG4Cv0BGw3i/wpWR8Abetrgp
D1fUexRPgR7j8wKqUBSr0GIYb2fx3gk9Nbzeay/0LH/qNX6B3Vmt11YHpJFMN7U3gFBFkYJjkCYB
Cvd/bn+TBMd4merVxoLJg6VpGPAsvwdgGQN5JuPNYFMSWxvEUpoM8vq23bg8/H9IdX4HbEHxs1g1
vBRrF6KOwZi581Je+/5jFt/65swdmEtoi0IqbQTGcSiL73IDCaxwpzk5xKKFg6WCIel1c57DaxIS
XdmRbpMhHvmVLzIloF/GtYPYcd0HOwSGiH2ZFSKEzYeF7EseZ5sVP9Tm2ie+2hU0wwqCf/iiD7jR
HRkpo9BAZs4PeIXW8DMn/1csjwX2LKQ9dMRQ7yI2muj+GJ8X9BvMb4+xPR+K3ZJBrXuyRcJ7eovs
R+4tck5UKoLYgP2oAPhLjIl2NMjZl1W1b/xy+6MAQ0M+mGIf40wQTe4Z/2+0B9YtxttWnn7nvXh4
iui7HzH79CmtaRCxgl+h27mAPOMZoEPUj0ENfHP7/+kyHO9muHyaHonYvFrY9CaaBj/LVR9D3fKo
Q7HeSAZQDx7f9ReUJtpSPWHAJmRoZ+E+ZCnA1Jz2m/IPNK4nm8TE6/k7voP1YRSF2y6jotsGhJvF
xG/8I4xOIluPh/SwBc9BH9WX8/FjwEdw/VeYSK/LMM+WqKQ4S+umRnl1sLZ5nKwDz6AbK7lFAKUa
kI2fafdvq9WEZEbBMVwVc94yh9bI+pSIh1ejXWrNG4/NaMqgWRzOziZj8IwFg1hxxPEbUdHNBqMN
W9gzjHiZsUXQuiVmqzg1biSCl1mGw+gQLGaF/QRmFlg1/ZI6D/BgvmcowZ/VyRyWvA7vQJe2mJ6p
O+vPb9AyBXr3HSEPz1dvHAo8bzBL/HjPNohI8/6pd2CvR7jb/TimTGMPO4xxJQp+L1GXhA/bs8V2
G/iHIZ3T7OUj71sqbEzdZaFiVQBfQMw6NMvs4ld2J8jQ2am+kxB5ECvXcTNh5+DIK9CQFeKgVbvC
/zdtmfj7B0bxQa2a4Iq1eoTe11U65lWUnxEx8g5BoF21xoni/cG1F2RfheE9Vket7LebhGqCZfBL
NUV+aCY36ptbKD14MgTV0fTZxgSzf93QcnuJiYrBTlOjgWz5AwgRpG7W2Tho4xwQ1j2n+XB2CDO5
webNGSF+/gJAuT65kRUZ0fPvWKLVYINsfs4SREbfGYaGd9Kf7qx6w3M1kK36xS2NgaCpgUEghcv5
NURTqEJSpJ2MDYFI2UumBE1y2hQgqrgSE46LW5GhU4eL3Jh4neH00Ll6jZsKvm2IWpkx6sCSRy2O
DIFDLLg2QVbPVU0WSybaX//o0za4RsFw/J34/hGpvSSYNqdVaIdlSgSVTr6kpEZfEOyhNJowI1wm
CDRmHKT5kS+84eY9F4Sqc+8UUiY5Rc2fYZ2d6HjW8gXkbO2R0zDo3AiJv/BRtNjmPp7QrZXmRXGv
0WF51Pc+QQyuoU+zY6AN/QbcftBEU157D+0fxU0SEERYILQIY0FAQho+8rhS1B52aUDuhx0cdXOP
ZqpPFHUzoFqoVL7ckJH8qDznWCFdFzVo2mayOMIgZN40x2Gwn0gl5nOPJIpydmBWnt7nqZaa3k8w
xuvflP5P9IkJu0PFrC7JpWHvQTAyouRViHD1W4l4sb0Df+bmBhqjG4yU6l3pdttufTF45J1F3ss6
5cGoD5jrFSlReLhFPBExiaBD4DUdUsXqQNwQN+g1j7ETlLSkHj8PSw3WCoL9wmGaNwGyodHN6i4T
vqyEgxWwUtcQY8ml0DsB0bmYLHgTZnDsCjX+d1lLtjwQXbWaDwVsBTP6LTrETuMikvBoP7+P4CPw
QnfiO2FmZf3d7wGSVbErOcmx556NEox/RvxUrtW2PvI97hOYZEDUaKzPFCO2E6CA6/Y5Lw8MKLSm
KR9XC8ula1fgjX9yy+rpvdRafX7iDu049PDKHFL3YZWLzU7vLQCf38XvOEyhGKUPgUjEfO5KhW/Y
PVoOIjimGrQsDVKz0FIvaZ/y6cZq84/d3e/C1UBLB0iP1KqwI3Z73lLqOBnlN/XSWHpyugoi2B7G
9oORfoqgdb0pDmhv6tXGQSKX7UHsslyGvLLGK0xaByasW5Oa9v/beoJ/IIbvm6NV741juo4CqHZ6
JWUSrSyw/CHkxen2E7D9NP3sO4Sgho4OxZHu+8K8prcrHcGGQXE0/TjnlWPkf/yXpwxvjFoAhagB
mxqmwOB01Nka8CdT49Bijl0o7BcUj1avqJ5GxTJ7+0I1Umxb6zv6w9DbmogPmDcyHRQv/lG/djii
mdo9L+dcnN3FRa1XGjUqFXqzuyC7IW7R7RQV5aQ8m709Kp3xjQwJ+/rZ0UbvZ7KrhXDV44jnEko6
bZ3vUtVMowsaHcIkfH75zOm5UoU9aQEOV7CSEfDWXJlYzsPk468EwQcJ3A4+iSn4InanvgV38OsE
egsnBx7rd17z2sXZ7sSMDu14QfJWFCZzPQh2JPQBgTqZNM9Hbi343TV2Ol9hPjsI1rR6kg2UXhvR
UpqoFPcHFI5O7/nMPbMLz0E884XnRudPgZuZlsRLQoaw16Qi71HS8LdQ/tRFBh3L43/Ul4n+7RvW
1DijDs6KisiqJj1LHFI1pHcefxUg15obe8bYpnlz2xlW4MoxkUilcuetwRDJpuCw26uxnJSUinF6
n68FOzLYajY6MxJxev5rusdLlTmH5sEf4wgHmeYGZNCUqcihDbfc9AOoFV6QiGif46IwmgBYkiNd
e3EAQ+t1Mry7M4r47zX0GLqPGfdOqvUt53y9/6Vx1n31ooC/u/3uI+BuL4Ck8+u5kBlvXKm0SIqN
FPoz0JUHfRYbGJEv0F0NTbNiGIlTIQUmwzrZUAF0+zKDDgxD3CAcb2cThqJtF1OFOz2Xx5YvfLx8
CzkUUyenrHKcuRUoJybQXAUUJsFVQUazZdIlbsJOhIut+U9IIki25evCQ7IS4Ooh1bcitrsv0y63
vinAMQS5kCHQiRsSYLldQLx0Qkppn94WoYhGA7eZdPOvZPQtBADZ7juKtfEzKmQD+a8NUNImf7Iw
9xPEybxY/7jp5ZapJj54QAtuj5blF80vfxp1J1dZ/qtMxJJJnABRwu+tjPBiategr2v16PrZN0ou
vPhbzshiscxlxPDjQydC1KqJcxZCg31Q7QUyd7B3+H8W4KZypaeCwqrWy8S9ijrJd7bfad9ZFNG7
SfBFlGqQ8DL9a9qdhd13cVZ3Lvmh6mGYpfpodk2QIqBQDjdS6MWINo/Z98Lqh3sFLkA7eax03oA+
qdwparC6x787PnTTxHpo4aqDmErBav1Sc53PvinmUIICed8AOrzk/uzuGZi6kkF4hSPpee5xp/Vq
V/7g4GMmPenzPpfQz6O5Z6O7efV64MoRLRqhGBWQ4gFSWIquqtGY5WtE8nVh2x/KvBrpH2Kx+yxO
bB3+ZuFd0V9iFGnrrZXXlqHblcpqV1KzElCTfe5zYXfYtnpawhEVc5E79U3igRoGwASUon8fpUo1
Tfep9KVTxU1xdZcHWB4TGXtHCic4GoAZBD3pFrU8dB35uHVgyZSm7y8EgwsQDZNaBLDjnPklVZeK
8fz88S1DyLxh3C0J3jkufu8nPMMtyNGZJ9mnALAIlQLMHq+Hvn014WsqbhWvWlitYGCJNTUGpRBp
cnTvRlAcVS+s8pMhwfHVrE2KxwjNpSwGDuGPszWl3zZTilSN+blc13+ifwubprAtB18jiOJN5ymN
hcSFOhO5MU3WaU2pTH8M4hvFy5mYTsypWwBE6J6OQqjyOoswyOoZBQzbSoI7MVg+IDtwik55vr7v
7hFitHoS2vIiA0ZaOk8ToYSdqjlm6hpMeyKjaLqHSHxjJaobJTQoXYRW9Ks/lxz04s6HNo8BFV9P
RYuykSk4b3cMM5ixng9Cftz7INoh5UcWO2Sj5HZt4Np1rfPhDMDjssyqqgtalbdCmQlYOdZZItDa
ZfAvjIS4ktnwjiLxlInR5Ul/hNxVhYG+T1sjf/mwdiAUjViK3nwVMlrHd2eqs0kisZZsuUvEIBw6
Qk/8XjkDUkadJPLbs9hxAcIUrQ5pYsOkBUmNtzZaMbhAfUWo0E4DqHvRr+qMrpEr1L4iiwZ0fhpq
fxE0S1W6MYYeus1B7qZaQR050weUjFEwQW7H8nMBgFNWZ0vLwgsF4QNj7IeXAWkD31lTqFD919GF
sBKDEZofssrZuH5sJiIBmdsdzFvGkVRHHUJxWr6hYcWz7ZDIJtmO/IeNO0cNQ8Kwlxb6V7WXT1rL
pciuuypBlGBszvHiKB3eCZU7mwILJJLP49gjRItauH9CsmP6+C+ofHiQHDuAsV7oqNTxk8NHKevs
NVtHf7KIKMexYYijPxIFGFG089UE0BCVwEQ0gZkn2QdS9Evkm+AO8TmWCjRH2FCYjdYaJ0mdsVRW
82V7vXdupuxaqqvfXzrdZx2igiDl8D1CGzr9e6IjmYK3V798W5Wpod8LzlI6VSbreUkk0sncAquI
tFQ6v5Zwid5zgGZhgcjxcq+bvmT6vZSQzxFfSEA2Qmei8Cq6BPiT0rYeEuMEu6GGHL+h1LTprwdI
QN/rdLJm7vUk00aIcLnOMRv+A75oISgGqtuoAzqCpdDSfo0BzVN1ApiJoUwz6qunKhglnjtOKc8Q
0nKQXMmbTOg3dv76bwSLxfICtxgfWx/5BPs6eWDUSz0GrvjwyY2Ilk3+8Or0zizAKEOCElF0ncdy
28FCxLggyzxsWD2w4WznQkHDJnGXxqtU/w4s8qZJUVz8B1woQhUgvW1IG/li1Qdwd9CuzV+HE2xs
0u1HB/3JGM9OJwTIZPTNRbDWyt7QWHLwvNOs/Q5g7YXPbJw0/HAYFeWP7nnZto8oimCIs9mzp/Ud
7h8lb1YduP7AKTDfp9IBPjRDpMH8D8gU5kIc7ueUOlOMmVgI9VMMFtRbw43782vIS4ZTNBGTSmtL
MaiCRMdOCaPPn5LP5WtMrUzNgWVpWKB9w4AAg1k3s+0PmHNmwMxVWD2Mf7x5uF9Rlgy1b6FcDoBV
C2xR+9pHpC93hw6S41dRsDmcaEeWbJ/D/G96T2SXGgiwWzGxWDnwtfZMMh08q5q9zhlvujg6NXrQ
0+1Z9gPbxs3IBW09m/WBUtTzBEe3YfGvb71WGya4K0mGYuSOuH5I/eE+V/8A+hq4Gebe4hoZRPFw
ynkTfqmgd3Lo6uXDhE3hisyfBUwnmOVWC1vOj8PhqaMivBMGoQWknRWYXCbZdNY7oKxJ2/Djg1Hv
STFFm0PEm1Cs+fVUhfSi0GN+dbcCb1mXqAANF8z8VRuabzw+x5+R4+qRozn22TNDeL1T38x29cuK
D7TwXqOwCdeASJCcXsddPH0k0Au+HIsfHLP4BD4xjsbmoFfoA+bNljITaF+qKmcIP+7wsWBbScZA
/Cc8Z2+oTXYGjgk5UxrjNyJV+d/n1CO+vXhXG4VtXw/SvWqJvtSb7bv62IREmGwnHQizZ1w+LILK
R1kZAkaBi8RL+J+SfkWzOm658q6ai1cF5+jfLBQz4lStjFT1G8WZafuU4byGwXT+fFcb/jVKa2wV
lzdszDBo2O8/LD6UfCn2oZVN0aF4G0ANzxh0i6GMDNl4l+dutbz9no/Nva9yVm0ggMU0dsOVVKYy
/Te+y0CpI3ZbKfv0WlYXYdA6GZPy3cKzcmy3nH9zYxXrDXcngnO7TmtBbrVXNuYmXKxpCIoE9Po/
6HUqUyJIU28NAMJ05NLbgywVCMRjQ6C4rlnNak4lY5v7i2tU20f2l42622XPMo2+8HXM2alA/i5S
w7OkNzDLtddlhJ3G8vWOEkC5CWWCIY0vPwS8iEVxm8kHm3vuABGETPCJnPC7iqJ2JVIhUwgECPf4
b0OAGO9/lZlbbRb7HPvqPHfvW+XZvWyNu+6lkBUW5DtnTH2OcZBbDvSCDGfi+0Q2RVw5okr1DgEX
9LaEYprMHzAXPYRtw00AT0E/tY+uFDf/oXJKlTg/V4JUjYS8uHdxahU+3APHXRQuEhDsIwr6+WkX
hpgollNuA+KUzA5ezldOuabTLpHZumKuaH+ii8gYk01YNXfO1ieMTh9EsE5kzjX2BaXEI8rKDoZb
ptrPQWHajqYK3hKWvkvDa5xbJjGv+TC2BtN2trKrWYvjYYFH/+XGb87ZKUJueFvvQhSaeP7t5LSg
XXioRqqVF7wBWpuG5AlOnDkfbGuEafi6uIFVoRkkUEDQmwKbLDpiwAPCMi6fN1cTHiqOz8Y6Xdp1
hIc1JRc8MheoXat153XoFiG5rgQBf/zg+3XCJsee8EbIjwZTErB7tIlinhxIWcpkHfRq7q0y/agr
zFzlF6UE2zmy+o4JvCWfMo8YJfYwf5WqkFcJl1FvJPYMyg7jeEvi3utEkN+hm8uJ58RlutOa3Y9+
0nEipchnS4xYTbEdGKcWyGmOypsIxTbaIEI3YyWKdpiXj3HH5NHc4J5UPteVWKKqbDgFNwpZ4yIy
YbwAdBwxzYg+OE0eT3zXHpBsUEz7ji0r8XQqEV0WQAaRjcTe+3JuFMaNeYJALkWIG5oEcD7pfaTK
JtKk/54VlF+sRt8hBdXHmp4efrd5r6ePW7LmoSs3FxdeYTbCd80barYk7apD2f06Ky/n77bHDbSk
bzYUmXuuCOwNzn6fdiUUxC0AwsbYS6EBos0DRda3heWcKcBsa2Jj9ZzvfXNpVmv5aELUWLBoC83L
5bOYm6rMml05deiqMz0WMA7N7QF4/1dUQU/yDrGB8KhdCcGMqtydSxDs+LmPfYE1255WGIIvHUge
dPiQfVkPUl3WE1TXbINjLb2BpfappZ7ByFbqLhzerBj0TMHBRDG2R3zfVIKO0MxSxxrRhqACC+bn
JyXBYBFlPSkT+h7AA7Dtx3hLDUDwNkAn577NwfyJa0dUdxgEvejsVV0+yKrojcnTr3AlyC75FAm+
/yzwHe9580WPv+T9WxbXRsqf3XdcJlmrc2m6lzmo4v3auXzR4lDw3hDZnB4ZsoIBZ9zdVP5PtI1X
jkd9mOaeV5nTX86N5DYsY9/mQDY8QygA3mXOuAQcCOUy6PvudVD8CvOtDi4qz2+yT0rzQFo+P1fS
JKr8QXe9vfRYdJ6i+HwhBO8uOK52iDsuAwG+s7Y9UJSCex/DR6netzsiaU96xiDaks6+oQB2x7Ly
RF7RE5FGsVC3nqcpqmJYHo2jBYxQLCtb0LAMKXTe/1eFl+6RSlyAD6Q4fqIRljiNh003x6gBYqq0
GqRKn4FPBXpTxhSHPYt5JaNac4nLzsTilRyi9f2KsEQwDeo9Mf0i7VrQwxWzFeyZLUe+BhIM0Hux
t+Yj1n0PoAVTJLZA0HGdDMHQqZhTqAAfvZEz/LZiPOe9HB45ggxxAaHNOGYfzearEOC0xHs9v4EX
xSd5KMYgcRR/0ntFgJk0FjaKLjhFm2B70pyD9ln24Uzkc9zUZFLy7X0lGNE6Ae1h4EfLRHTPc3gb
OAb3k0YhFwQ8paW0foi6wQL11gqGq0Q7vXWNP7I1G6C7cGrI/FFuTrThZMIlZUW6kIWhbF7jSPAQ
yn97BtQdrqHTNy31dgAWIiNqaSTgvC0jEfwuPPh8YKWyOHTDUIuxNREVRu5nofN16lEaByZHwIPz
1VjEIXZyw6tUf+QZYIK4H1SaVCk0kTpNLtSyYvPNPV9r/SA8YpJylm9EOHTtDFIn17JGnR/aP2HO
FqtNd85VPhKRCRdJuPeN8aHxMmqDl0z1pEcX/ah75W87EZyM/emCETQZ62kHPIiF2bgXrwVaZri6
5qoqkasmaScI96nZRCa5YJhXVhuf0caSnPMthyI0eFVBFjHA/jzCljfxfA4i/8koKajejFHPxEci
NAEWce8KUYqvXUEUwa6sV4vn0V4E631lUg3odJS+WsXhgCyi16LDj+HXe6cccEeSzBS/np/kYjdN
59uB2WwzwDFp5WBr31rerBmuPmlSZD/629h4se2QPI1JpUYlxtHNwL+OoE/0nNM+aQHI/rYMrAex
Vv2avSR2/C2pp3maQDPgOkU743j8miWoA9DFP9iGv+r9tnaBqriqTrFJQ86Occ52FjfJYze7g2hs
E4ENUhs/EX/sq0wz37NudXEgwN0xiCDbWM5XfL7L7E9Z06ErqXVLEWdxxDRw9OVvtzDgQz5x88Dc
3CKCIszL1E+WMfW85rhErqOxdRsTKWEiCDge8q/Ax/81GsFPIU+G+GKMnp9MTTt5QctP3CpBsOCA
g6wyoIY986B9NR3UqMuDFjWOZJUsU/5TYW7iZ8qEbTxend498hmmQIW52j49bjzalpu1ZpaXe+HY
5YYPvcNOkXsWHbEy4ccxHZJjy7xQD5YiFKUCplvJHR08rD6z+VEpAZwiPcCJSDNeEpbbg9JJ/j3Q
3xHLGVBpMI9tGSqUaV/ha3uRyFHs+FkqTZeLkKKOlexgss7hLAXA3OHPQI2y6o9iFk3rqR7F5ofH
0LQezTrlve8ypnp+8+4NzrzXSOzlT4JrvmOOH73qANLbSkcD56MrufLfcO8GPtiXSXGgUxUNC8p9
XdlHyXYryMKIjJfEyWLh+q0t+t7VHJtnhMQmwVGS/Kxr5kJlHPfV3YEl6L4n04ZRlppMIDHBZktE
vYtKM6Z61A/MFK7IBm23AzdxVkWQ91GpIlOKfXR2wtDBO4GXCBcERqqwmcYUpSb1w6+PbzpoNq8u
Julkacei+IEdzGEox3PzMFLoFL5lOTyFK1yTMKZ0yVNkG0mxT5J95smEO8a5Ll1Q3mPAD3cLdw70
4rTa7k4lHS0ps/dxzHDvC7dCADIy5+pMOVwc/eDUaOVVPQHGZNp0P+nWfW2pLwVuerzUoL9x8a6O
Bmp5i5YImh+5JmG6gSXkCJmbSNi/TNh42z9NICwyyHp3YFfjpDmHS4kTak9Bi/PyckHOY6v8Suqs
R1fey8F5CPyyqTVB0h6aCFbhluI6Ilgey2t72ySy/PWlle8rAGjryohvxGNq++kokjpsGHcDtb8p
BxKJ+otLe+tECHLkUtsuBiSihTwfoJkZg5mexYnGXHGPYgvKfHny6JVB2Pbwor5xzSjKbd4xybIy
2WJRnD6Kvh+stS/Yfi65Q4H6+x5C2na7TWZbaLw2G5UKNXvSGE0prJ3wzp/rQeNcHBI6UdAOAsbm
pUVDsvXkQ90XudadioSG+10AP0VFB8G7GBZQvD+0VC4sstFuPtUeVAqCiaYKAvoWwxgYsfOCZj+x
l1EJUjUSJlketDF2wh9+aIrwtQjsKn2QR9NgFIvcKmLaX6tyhzSUy7nAhvjflo47FcRi+HKZOIj9
uGB+XNeaQ1BCWax8LvNoJwVx5zosbyP9S63KboDSfgVew3U4oOkdsKmW7GSNahxSpaEoihn2uH6M
lox40rNlaFsjHfXlv2BbqYt+1ycj6gu8rr9/I0dyF2ECdVdN3+711jznc7WknvTjvPgDejiNtCmY
jkkYyKZQgPYvt7cIn9SeXy+vuGdtbnpO9kMaD46TnoXRM8PgAGUlbov/NBvbjagvMLKbWjzemxHS
bO+VHBHdNVMRqKYCfg+qdPt20mAkdLKm7gxcyotbiVVUnMOzCnAMrpJStpPh8CQSFVSoUtJxNyxD
LXh4HEOVpSkA9LGPq8xpQuFDK6cXBT2hBWmEqGXdPd6cMXnw98046clmu1oB7hRyOTlCozoYnT92
QULO4hBrNHtDenNxK7Gkt9h5rIaP/QHAyqorJeMPxprs+6l0/nW7VVQV1z5UqJqV8Y4dO0qvNU19
B4E/U167PQToLhw1zEXFfg4lnTaVH6jkLjGnwS909e8BXVK/0KCibyD6hTj68hJfn0s4D3CHnChz
LHjjX+Gs6bujgmOlsPEBjtE24TyFvAMRMfYntGt0vvBABTPjLFxQMNYFLJrXhCvP4ZnxpzE+loZw
R0ufUVjXYwNx4Wd92/+uqwYb6wux3BHT+z0mCN4vc+REJDPo1Yd+WOpbEe6D8ghgFVZ8tJ/61txG
wIiqZXyhUNbCe39KYIteZY6WRRhsuc9QAWcsB6X6QOmsYTJPFoo5Qkl2LoDPlBw+P3UCIyrIBdsq
NBMsolkNYLDbdW+1fc9h3XqTOBXzS+T4X4evwT7zmeQ2oDNHejnS3Uy8tsMv3F1JlGXCyrLMA7GE
IaWahPY/ktnp3RFmBEfbLLggbrYwsrDQ86JxUCUnIqIY35moolGMBHS5xuCm6HlZ7lT8Y1jnbdyN
Q8QRd1Ph+15+xuUi269cxtudt/i3yi30Wl5BcQ8Y40fR1yG3ugq747ZyjPIR/IDbyjsGJPv3q/aL
fs+gIy9pkJfkMMGgnmAtFyZlqeXrmN2opIunK55pmy4l78poeehWVDgGZUF2FwU9DmTDJXOUeMM+
jsR5lyLN1NgdYY8rn3i0heAci5jmAupCEJdZzeFppDQtSUgD6tcgRSBeC09/8zXV3T8996tWvkY3
Z2uXaAbZa7P/0EiHnRnQUc2Jkd+DhykZW2MUwnXWow3Cg+Hdv1mVrVzyr1E0OfaDLH2dbneHlobT
Q/1uoQ5ik3HXIKJcvrKBUEcGR0ouRLJNZpV/2R10Eky/45ilX8uKhkdir6xSRzaiSMTWBe3mpy0H
xeqh/lbmlwKT3+GmBQwEhYXD0XOdLtqRjxSXfoCBuqGV+74Xzze7VUeO7Qv8SyULHz1KQJ2nrrAT
GQA8IXFrx6A8NbCYsHrwqfo9IjPAzf0NwxNK/fOALINUwMFNO5x0Pk0yk5/Pt+l7OWOvuOlUlKn7
ytBL8HiIC5gzr8VVkjTUzLWEDy5QupfDfh2OCwpbKKpCZPOoX8tSum4ior19m0b0O8/4RHYVvVZu
3YJ/E9UnuFh9/QE++pts1ENPyHOQIubC39Rzp2IOihN3cmNyCo1pNvEzuuAQLgu0j8Ao7jJgtWFn
1TNdRkc4YIbXPlTWcVQNpIDvfjzbsq0s5t8tf7LJu/Ws7J6kkmh4i2LUykFYM85T+yqCllIQT5pj
SKIfY94gCmoO/Hwc71nllaBGfnY096Mbn+PGAXOAT7Ci2C8apXnqRaXg/4YI1L08Kwlbj8mtgZn4
OeXv50YyMJRi3F1+y8VHHor9GyXr+c0Czwo+TMq44qgcZZAsfrFd19Fomzar8qJXty+w7wLeGSPs
P9BEPVUGWylBsOu9ByFqtl22nUG2KNziKOOTuejtqqfS62G2ipN53tMnADgE24PEh9ZD18T3QF4q
DvWTThkkytGndrYbc4XWxvAqgdYHZKFqfjqLkedcpx6AGl4U2jRFLnh1gqxjA73ifMjz4/3PpbtP
vDMscD6H/0k7iFl8879Qj+Id68bm2AhQq5lpcJ7p5H5E5WYKZEGE4FcIzVe06ozq365kPCEOeFGu
Hx2Gtun7NZp8RHhi7ulIeiW/f83F31bIq6gvqSawpvun//aVygb4zbUIfEupRmqv8vBFInkgMftk
2yMIkRN8A9J8e7azBPBeDhXs05JoqecQWEL3afMYlaoN1iT3Mwnbr1xgg6r7Jc4YRjTw86wwSZ6m
1c7GzR6SivnkXtxOW6EFeqyUtL/C3osSRCseRHc1Pt4asv9SgWTiHTBwbEplFdlhkNvT/kj9nww2
AheVzy6k7SO2J14WtZzALTwcxc9PxcFAE9qbZvWRtCEYhTefsw/CDUprIQFU4XSUtVTkLJ1HW/3J
ttZKnakk3rWrdI5vYoFSHxLwKawkQOpwljh3GQEpC4hrXw2nU+e79fE6BBssbwAe8BipPio16vdk
oVKn2WbEFZ4ZKC8t/1Ngje2Cp5sMuK6lLi3NKFmLlnDA+BIIRJ2FAUlZb82sC3+ewgWj43FzaLjP
A/1b5pwjOkSYI1X7ghUIXtHvOXc+KsbpdtExrVjCBvTgKgpOG2q0t/8ooxPUBHu2EH2Mpv8enbXU
1grhL2qRFczsn1T+K8UvHx1VIrD2buqXrREgNklgvntnJ/7fE0yKiA9KgrGB4vgORuhHJFtYtm6q
jXiVnGWJaoaZtL2zlO38fr3E+b+G9wsghehqBDamMUAxdc8MDssb3dcjypWx4/YiiiqmnBM4nd/q
9nEtLitchSUHDhXK4rWE0Ggc3WVGFHGuZQjKrUSvbvzk4461kTMiTeTyU2w6YQtcHHUuokBia5aR
HAO3HTNMtk+TaHvMh3Fd7X+84FIA9Gdsx6+PW/yqgX5N3iB7jj3k6t/wKV2+FhfzV71VgV85Vgig
3uN7dnZ2DoE3w4LlPBoc6NmVSnA9RzrKZE9qiLKNapK3AeVqnYWZLfXaNYL/nRM11lRSrA/yCJNr
vYpI7/45yJdg4XcRCEuu1RmfMkPgZ089QQ3fym1wr2OEV+3M36l8wewtO008jcYzKWx0BinoyETo
NfCCB3EQj89bqz2tBOrWaZO34OdTsiLtTI5colWpul4C1WXylekEfEO32kj41EmLgOLcU+LUpwJx
6Fo8iEZn4pcYe8D2+1Ec/hfMCDcW4bPyIbmfGNHc37L/pfCUGzawlUn48uXPjw6xoMw2ycU+gZly
iR2p5YlhMIPWd2gWc9ofzgEEt+b10CgRVoTFdqDVJSSyrvOQDQV41ji1RVDdhGlKQySfFOzPSN9A
nSkg36ubSx8mEShkWf9k6V30MSrFe+hGQcAduFP4Oy39L+FcwOy7IsjWz/ZDbMlvnlJKtMF5o5vo
HtXzhgH2JfCjHW5ZP05mc4IPoQHNR1Of5zhjd96+szFfksLHja4Mwi5p8lIL3+Kvri+Ta5dk9sLZ
ocPGr/V1wHh/TsjZNJcmIkLMNggXhn+ARNGu/4cxp8mL2kwpQvqMTxUhmlqjJ2eqj+atlqO3AFaG
MM3ckTquTAVFf4BIfGd+rb/XftLEfOkdHwe/bjHqlKM0mPRaZvFJ2stlEgTSpMWVIS06OPzbMSoD
1zyhwspoZ3WUW/hRS1sj4fEmmCg+Ah7re4nDPHBPY57W5bHjxCOWHr9ffn0Rv015vX4XX8vBbncU
P46mDG/xF0LsVumPd4wgKBSCbHVwMAOeD2cy5P7/v2oZr+JwPeX039/oiV6uYWqfgmacFYnV0ByL
yRdgmXoEY8D+IEJMLCxwnF+TvY6FDpiD5uQoFqFeRZEg8EyllV+nJdMQVh8Rem2pLfg1F1lZSnhw
41SugLvJ5q2DKBKm6QZhGGrAU4sVzf2RIC3A2pZFJei0qMP2i0qOOu6ITN3AlfFNg8xOs6s5j3s5
6CYe2qXSlDm0SBirq8q0/8ruYD+1b+5b0ZbHtR0wE+10uR5IFTmuRBdCouwIr6CegHHxhV/Nr15o
c0e3/I7KPfRMDC6u57tsAmZj1r9mao5r0KsIwNuBGMKO40kfJIW9K0z3mkth6TAk5CUTC1BNMXxs
U6S0HIy2NyILCWNp2CmpQS5wUfO1xFvhbfzUqFZ0Q2HzYwht2ilZU4Vd1L9UBAEVdK5Ztbqneggk
299WFQklKQjnMWUEEJKF/TtYMFkJYFxmHVdzBuScg2uDkvU46yZNTMp/IbsyyLmSydgTeg/kciSa
LKq+WeqH7azSJefGFdXdav2laqLlXCO7kRvirm7zQyq27HYhFwZAUj21Q2uC1PxRQlkmFpE3Kjhe
6t9a3TJA3Jz+Ez3grV/+V92Z3hbGrJCLpxrRN4iXWWyDqbG174LU3s2nH9bsLTdN3FbkjOWioSnc
ZxhUD28IkHoRtpUR6H8pv1TBJlI7Y/Jk/NMxesnTDWk27lfnd1m+yfkwHO2+fjOm2JeCKWDB5/2n
RVSCu9BQ8KwILHjKn5H0nGK/CbOYh5KOr/KYUhVZdVZ72x2KzTmcs63m0y0b7cnSmChc5+MycjEe
KDer8y4po4t0sE5LflgtxHAgCHm6BbHofpNvt9BIyPnzySW+ZVtrEF0s36WHDiIOcS6nETGOoXHq
77HomXppmI/tcw5tAhJ8YSK6b7UZ2nmfueRlwsE1ecC1nFB6Tka1rsd0BF9p6s+HWRxkWyKdqSCc
QXjSMWgPbycFYEvStcHxwigZenRGGrL76EOeBchT8GM6JroDxROkx5B8B+/u4KxhF635YRjq9R1I
qXXmRut1Ljuao6ThT/lmTAJTGnooBK5hotKs/7pMhCGy/k0+arwTrOUB2ppsj91H6ltymNIXu6uC
V6DyXGQDB6wRUxiCsNKSTWY9TIRY1Z2r9O8cQ5Unm6TG/Hdj0BTM0tnuGG/jQkQH8vg/mTY0pZkl
2wxdyt7TfOKK39opZR+hotVV+yJsct98NHFmj/1dp/oIS/aXHw26X1qwPSTyo1w/Cp36m8fivPCv
bjCEeBA5a9nKwnCIDb5feFv6QRed+Xt7gkmjtfeBG+PbzpEXLY+PKWc8V0eWSAuGJIpHNj4zA41s
QJPp3vTvizSmtRPUgDkEHn9hB0oeZ26FXnNFQzgPFg2bXM47ZXGz7mtozV9pD7u8brlDZmEAXyFy
ZpW8IkYmwlSNrqMqSBQUxb8Wgw70GPAyrZjQc7J20+J+cFl5QE28AOFBGOFOanW5wDWHKjVTYvw6
JPxVEBR/UlOMOfNG7tS70tA7hw45Zc8wqwAbts0jhm06Jbaqv486ysO+031jJgYSy7v1IDviG+WA
a+JIQzBFxA6X9xK/z4p+8WiE7IJblDJB7JXIRqZ8lbgLZ+hkHmghu7IWIHMBLZdObrsyn4Ab0WNg
DksuIwMIz+1y9Ll0jYg0gevflRve0e0W4N+puDLS1ngzV+7d4zcNtJHO7yNyyoW+NIY9Z3H5dicu
B3fiv02UwGK27x8fIJ82BUvSp2dLyRiJtu4bkXW+ZRzm3nQGGmPGs5r3sgfeOuLrepo80/F5MrwO
IQ1nQ+YIGQsmozBhH98HnWXXLBLmSj6j8JOSaP4nR8c3q4PP3fV4YNctYs52U1t4LzPoNIfRqZXY
I6QsduS9gL2mP/qVS8hwS99ZF+J29b5uAS0zrDV/Humy3BJXoSl3Qx1qlhl+a1MRNzjVKOF5Uijk
h1CDmzxFA/VyEn4muLXnjvSZsvY5940O6o36Rq6i0ZwnCpgkw6Kd90ZaZnHs2FGMx9PCvV6GXykh
TFEY+rheEErYp40Pvh67z9nhkDCb0VOlfyfeJzMfB+Hmv4QTu/oC7ZKt4COvo5c3S2ZD0xORiHFn
mEdogbS48jfkxHco/n5Tc9+vgZb+71NgppsQXvLKYwkKXETd6h5oj0zTMkuQ1v2oEPaLSJG5J5N6
j5eTv5WFOKu3mlsExS2S3y/7Ik+O5yTDlUZH7Id0nMuZASRQBmThuL2/i6N6d+dNxCpPTYKQrWOV
c5mWOT1hp3NRVPUeEJ/ClGrlaC3QQIAck9p+s90gR2Fg99NisngwJM7+JM+q2d1Qlg68R9NwLuix
IwNXWKb6w0hWKzPBLmlQh61CSIJkeVjgOyHgaw2tAud2fSSWaHeRDdqSq/FWjNDks6DI+7xFTf76
BGaSdCjKYHqnmODRvFvQYCnAWCdFFrjIyTCJ8yRLNlyBKuu8gRPQOewR/Ed3fukuCcnutAAuF8UO
Z43QTHUXq3zJa2SOTJ3F4EiR4g7vCD/Rt1LspDFr015YWc7/988JztiTqy2azyYjL5Mo/+vXKkFX
aJpoYA0DBtXcYvRVc5NPfna0tADQocHOcjMrdDVsZeprrSK0rkjPu60xw2AVDU+UFfX7C6lZP3z7
/TpEMfTq6gT92jQTBTTpwS1b4gOdKp4Ejw+L0wj4N3sRhjLiZGHMjLZJO8yogwo4PjLzYMimzuku
/Lr7qHZP2Jt85IWdAgNWlXPQnFfjTJY2bcATmoS77m/v3wEKac9FDeXEaiXWaD4yr65R1xleHeZj
bUl9RTv0uKgCw5Zqe1pL6tr83M4yI1sSc/Iq27A1dN8qtssgaMXVK81lSZ5VT6s5ixo/tbaabKXc
Vv+qunghUedPO6pZ+OsD4XJffqfB9ujFhD7fwKaJ+3b+dJmwqZSVOsq2hcPk7Cf+h5FVSh3q6LK9
2tda5a8kSAubbxf52zwJUkzN8KPSPZiE9ag1C8HKpfTGWsxIng7HBenL3g2BIhOovIib92ixSC0X
eCu1G/YYT80b4hKzj7jHJ00do4cLlqd2uwv8FnWJn4+0+DnLixWLxeCanVig2XXnm2XoK6nKFVLT
T0h8uwzYtMG8Gv2rMNWkIjxV4D/TrSFpm1//0yU4Zz3g380qsoluEfdpxcCzFcyywetcQIveene8
kjKOPK4aZ0g7WvIkjuPEf0PTuCHQ9hfRjX0r6Nc3scInzsnIyCtf+rKtDWsb7bgKnhSWsU4ttD1k
L/9eflaUMJq7wX42vGTZggZ6jHY2bJWiaqZxeS1cNEMzbzYmbYEqi25h3f9IngWX0R8ot5qWIYBY
66U2WvOSKejjwcmp6cXiDJRPcOB6FBHrVkyAiahPLMauD0RhdW+7bNNC7zh7Ym1FsWsaLVuytFul
dxTtNZu76ruyOBAaCyTYKkLP09VF3B0n6wZXlgyhr/igiaAFw1ZSurZHSRTPsuAHX3CBRTyQFapJ
M2H3Zm+mGnAztW78fkzq0eNz56ZgxbjftAMjddGM27dvrxGzA9tMDT2kgDNAVMzsaamJMnFFpGyV
UxPV4fcFGdwYNBGwGCJ5iVhvRsd/WthZd1De3qsqTjEQ/XRF/Un10ZFJDjXnpgl8JvoVhnv4Ap7w
pkkqfHYvqZ0AELaQhinKbAiYykmIUiagQ7Zyly/ehGelqsJtM71swlwAVMVWaxL/wKZ6KfJrukXd
mNH4p2tPQVR3ev4IEZZ+hj0OEF2q+8373xdKNGpLZ7zDSxsPOl+04f4LUTLpr0FGFfZinzqt3aQI
WYTFWQpLVipvTH+bI3DbAsJGr/8zyo9QcKxJT3BkjQkPGgYMVLtc/a2SFz8jZJNXUiGw1QBm7vB1
0Ky9lClHzc7SuyCbQYtr93wBsRSNnKnYQXcAAa3Y70tYRZcG/gCIGUJ9OPqbQrClcsVsM4xIP352
r7X2kmvs7JVfMyyE4pRusGjQuaocT9yqFM/YogpYxxWjCj3K2VKIxAj1tpfFc8VoHOnVji0mK9sv
ujJJaYf0xXUxPGifgG7imQxvZEpwFylvCQx7alDWD8zBFiszep0m4iGoDIc/4cclD4z79cbWUg0/
gbTfBYf3KDDB0HhihD/Fyr11R4qGmaO/CDNMl2leUBPC448nXiDYYwmf49q7q6fXJG6vV6ZBkfeY
LKOu1VubYFOU07ZZcoFLKJyn2axZyJiueplqZI1zWXmsZDyWZUeGkfMfDs3A8/JWywWVyPSzmET8
KozoG87b0eiwYEMsvc3bGKC3j5Tpxb20b4tVi5a7ULNHgJsq4VH823yoKgLofWzQMGMDMuboZPkY
xYCn+3VkXmv06Kn41WhHjDV7RReHy2WlkAcV407aidkWUHR/q0pOVLkczxL2Y0uxLN+ep1n7vYcI
jVQaBZyuJAQu0rZT3CTYdHUPLqYMxlStfPkNqpBy9vSBtoGsoRsJ/OBNFl3T2ac2Uqe5LKe4dNbY
/EK1w9ku4C8ocYgpwK9qdHtW7dqzAPiCn+baE72xGWa+4YbFNSpMwmf2/D7PZ2mUaL+xVismW7o8
TwIL1Vl3JIXegMS/fnEfsu4S/LPgqhBE9iRXQHPvNfVXZwNLMTkiwSZYYiNVeQNrGdm0KzM+Yv0+
hQzvjSNWyEg2UQK0VHS63+FqDQHVufu2zHFuJlOEBHc5+j5Ygh2TBreDOgOSitsuxz/Rz/M24OYf
cqhFI6Z1UvEHAeVblgrlRaJewHITU4+r5i/hj6KJmZXXhioW5EyOcv1SgeTJzMG9Q+XR3b9nAgGl
ZZJ3cVt7UDu8DRvFv9FPusQ6QmMDNotOLmgrbV/fYclbef2J9I6J8FaeBWQLfIzp0rEvCgRE2b5c
RxwViSTOcFfKSccu2YGsKi59USEE9wWBEnsJkktuZvsuqnVccJzSsgLfOBKaX7HhLuZu0dZriKG/
gLZaz9LMUsD7SWJZ9Mh+ZXlHcqmZ+Ep02t2JDiL0d+HzgNsIcITnOy/JCTMk0B71gFEMvDb5WrBn
n0dBkQilaCDSG923MZX0/BsqPh+HYy86LOO3ourJtqhuZMJQ3DIqcQczexp0XoweNdyqNO2K+EQA
B5OF9coMXspXyv1P6uWy3blGd8dcjhi/88PUrl5KRzWgPHNkCUwSAsnWz1+3y3wvynr2+on2mIIL
wEEaeDr8nA27FdEB6b/t8QBZtDqU+i0l5MSxRpWPssYp5Mtcqgh58wt+7G9NiwHVoAsHp4/0hs2g
ky3M4av3GUCmGlYGWRSKvGE2yzFaRSU54FFoVzZ3Sq/UE2QsBEkWmzNmuiu6DKZkyYSV3HCnY4Iw
hbBXv2jxoSvl+9ZWDRoeL2j7m9kVEZUp/itJAR0V2rMk4PXogYYDxUj1cuXdH5Bhsu2h7aDnep/x
qY71L1aZq64RISDV5v+6pCMpLN/vEjol1QBKu74GiChJdMs+2loeZTcBIge99OeYchJ2og2khbn0
UoV36oU/76m9+lakMG5ER8EDjK+VL1PhhkB+DrtmQUcL/gb7VpKzT9dpI2WedhvKb0EHnBFnHym/
2R05Sl01sB0/hdaEfWxjPgaOR9nG+p8QnmkA46DZrfTw29AwphTM2ghyXrAPJsHi40S60o0AaYg8
JjzoyAt3qxJs1xg+wpT14ou8pRwseT0uk+rcnG7e3a7cjXDOE+YYstgtIJqu9+A+lNtUZtg0T/J6
OffEV2nTCJ9Gjp0c+bTNfziZHFnWL39K1QGJ8SPSpbNXASQ9snhsbs9ngJbf9JsIBPRGK4VYFx2V
7ydmkaexL009gD+jVjoOjXVSD1/UE5J7PeobjaGyn7OO7U3pr7N9ko4kcdo7MvJ4FlYfMzKMoGec
+DFibT2mgp8hUm5lHD/Na1dL4UyNfrSVoHHQevVAvTRTd86dNSVaZP9csJ+sKeI2eypS0s5AEOvC
BaIr5bNBFvHe3oKBRQPn2ap8AyjNKmQBdv8+gXNOcWKqoUwAOwbyjtHiHEKzbdcYu3HtwXrrrN1+
QOa/C7auDl1tvKjMHB8sTAw4Y0JcL9rNj9YF3lM7EUfz6uJiZXiFod8X2fHY+snEYrS69VC2MnzE
HpkYhkpTOXdgeZLEP66Ua+BQpzTJgjMvLfoGvqEM4g4W4da7vHlocuPZG4iC3Wcz6WKJmsbu/M/s
lkIJAcQY2skqu2VyDAPppmYfG0l65rDVaLJgF64QWS3D9bNr4ZvWdMDbv5qwMZ4uQNpEVrbrBVfG
nPdwdpyuRS2v7E4/a5LK1UPKdREUZkstNioJACy6O4ARse8nFu+CqRYM47IEmjQPuHZiTmFmd0yV
Qt8aTPgUszI4CHX18e4oN/B4s+zEFGyYqqsvry3i324jY7f7rLUwoY8ogUF/dpcN06FZG2KbAG7K
srzB/IFxjt0NsqOma9vpWFTwK9+GKXp3cw+RtCnCKW7IfGGG54Gn0hFk3b4wGaMjp4taXDOmewzJ
8hV8hEEaKLKX0MvobDI05DLW9WPImG8Rs2GYXCMPeVjfNl2SAaq26LwBQ2v3HHXqbBE8JEGjUQQO
gmhp89rf3FmxgVfoFJbEQiWTTtBo2fyYfCrVhqFzw2/6QJ5liNZBs1s+vafkMwE35OXkDt8AWzok
qwKuj8YRETaJ3P1pt7lG6ed5+mRCnXJPS6BaTP5fMMpQGItvvc3z1cY7q/tK6MNEeXiPgb1xnULV
6EVfg+u44np5q6aKkCJZnXTETdWuLQEnv56m5paej/A1kBy943b8TVmuKZwBe7PrgrEUnX1kFNTR
EpCaiEc+IYy9XYLGn7zTnMUe4CJoMuza/5pCtTol/VHfY56bVgTgeFauF5DdStgW7CgDPjN7wmzz
lVV+PE3irvApNshkqRxtTwVmUEg8yLtxiUbj5QveZmYo4HbGM/1j+3i92LBR/X30ExxLyCtnQUVw
Cp5vVU8Lxn1a6m7Q4MZo0IQxEVl13USJDJM8CaydvPOdRna3o80yTPTXxrW3i4jBDf7qbj+q22L6
XpG66FgWJ+wZi//DmJ05yzDZzDHmQzWNp8SX4fjaAqDylX8kCv59WEi0qvCoPWNa6PkhwF86iAQ5
Z0yKSREeiBv4P4QGX4IYAzzD5qSFUFh2gSOyRo/iU6mvTtzBd0kbZAlrjC+lPrr5lruJjaPPOG/k
zkRjbdGiuk38WHk/f9oFEyF4nveV7vTttqgmWRFDM49ycjA5l29N5ZI2Xo9zZv7rmQnXLRljlfmx
jC/l5ExdbAX8NRSzPkqxMM3YbKzf9yDfRWmDngOfM+ZiODfQ3vYRDhosXsKhhSwMh48Om4WZJ0dh
+dBtoOK3sGlYp/ukDVT3b03euLtmbQHEZ8uCiYll67GY65VJALK0YU87vgutHhnYR6E51OMLFJht
P5pNFdyIYYmNqY7/wI7+saHg3ZG+Jt32RBM1Cs0bV0xXUWX89lrpLg4ry8QTRL5Apg2tFbZd2HPB
czJo4/jtcU1Dhb67WpDa0zMCjiTWmJK/VNBZMJQfNkZe7+dwuO12hxLIZD6mBqIgAC+lJB+OpPxM
eb2ZDacIh5S3lVJN0Hm75FMENz/M6yAtvR4Tg44NqJBWAdokQuLq0Eh+yNDPISfxxQgNOFa0FQBq
TI56eD3Q2Bv5V5IqHtHPjWx6MBG6Rt87eSK4azExaE7jT9+8ASs9ms3xOToqyeHlGcyH06n2HAIQ
J1hscH9YwZ8ehUjM2pvrevLOhWIvGcDDJSEMde4BSjYcortEufZ8OttqhSEcY2+ZVELU4DKMowza
RFrZlDB0qq0ErYsiRsT7AKydBZxEydUc1oUp4AiHTPEjsMP0Q/a72UHcyI5uAJpa1ZqL6JpRkkb+
K4Vt4apnUa0dY2vpXfbEGImdnAM3KXynF7yjTnF21W38/ey2f/mz7K4ZnyqMnPMx0a4FeacPZK2q
eNwZnL2jfK9VCF2mX8PNfeAImko0OuhMNelWG1d0PJo6EXkJkGJnel6yemFNuGgD2CS2VATsdjpA
677lg2XIG7K97eViXQ9TtdOhhANB7jteXLBJGxwSsZOR//oItZkITaMjWOkBcX4/2Z6Zu7+azY4q
n33wgVP2ayPTx0i7zvPF5vMx2TkC67HXIIb18kHs9qGoWwFiOwYTyDwa+pR/mfkyxNRCOyMTGLDy
8/OI5LuS2ASAfE+b845ULnwawGA3hF1B+Y3/MXab/zbbDtj1GSMdn8BTma4xXHDF+pUk880LqQ3J
Be6fT075IpdV002HzR/g5/j1ypoPUHz1SoQD5g9Jwz/ucu5kkVDsWlDBY4kuMUAa/URQvjx+JL8s
nnLO11SoXKEDhBYVxuW2KX5O1/KAy776CLC+sJDm/HubsICY4eq1eA4Z64NpbqLpq2TH1ZlLItsI
qDdgX3yGejMu5KwjunacW/mC9ckSjjsg0G437rbskzN14SEeD/9TRcRoNxYP6G0b5VU1QZyqwMrR
XY/5/CYjy34zDly3g4NkoYUuAht/39D2AetQOYte8L0gHF+/83jEYxHdDh6jhk+ZEwuKsOhpQ1pW
iQLa9Tq0ZTAmiMFyBwTtRDwlmn0AxnwZx4mcqSWuB4ZEwWUp70tQkO1nkOcZB3EKDnpIDj386Dcx
kgj9i7m2guTEyszPnL6APj10XKERiPazXFzeGJNk5rZtiBDvbRbYWrAi+yaBFygk1Hl/O0AIvZ+V
NA/NxqcyohrvLZKSzDgRE03nr5uvs/C0NZx3rqpHhw9i+op4j33nSZo0Ipy5r8F8Lu5CFJQG6HY2
ZJfumUvV2OSpxxntotxnU3hRyqAklwhGRfAEFRTRI/2N5M+BGXDGMrnJT0+r5SJiaq/F7wMYSqvo
WwFDvj0DGZhWOSa0g/RiObAfaX/KrYaeGP9Qnq6RN/8BAH1tgIViEqTDawaYcUKOoIPU+UM3QKKo
LWRYnkEPvvlQ/bdxvABfKnPRVbFVkLDArUaLPmlf0jSFOUDKC1AMm1MHJlf59MeMLgJD7scymfWN
/Tr+2Gtr2wGIsDW6wXzghrcTMOkAl9HgqXlB21SJ1muUwYWIaHAlo3soIbAwSNKxpNHVIbMi7y07
9vSEesZ7cZonI/WNT8QxU2XT7BkOmDlhdoy4EHhVOaG7zbE6yw727fcwYgn/uAWwEeIbO0gqC5p2
/lGXbQyNwYzBm5AP/E5jaXla0Dxnzr6fpTkFCP2O5h/A5qxlngn2uYRGOW5l504mFr84P3sjXIgq
eyFn7+FngOkEh8AepKg+hZX6fx/DDf4dHszOz6nUEa8JponMvar9fY8hxNdvKBg7ZtSF3ZHcglJ7
uumeB5L//AFY0Nw4XuuMIyYPmS6c6Xa/gjlbzxS2TMVpCF8XLfXwWPJmoaS6S/C/lpID4ex09Wa3
j7u5pbyx3ZkA/sE3D5PtI3swNvwBRn+R93lnAHGcrpCEcA6sVbJcUap1uqfmadmhoV6i29ypM/ez
SEpViqkUowrnFnCjQiXsbH/ln8Fm0n9BKr524c2U1ThkbbkHq/SIlzvVWjyR06u7ETIExl8d2rcz
e6yJCZKa1MiXg1kZayco8xjFC+mthDDCs8uuKXJytAqJhB6HWFUfuXyB0vgLzaRh+c3dpvGjOZoq
G4uL0JPyGf4O1CIki+aUd8fpjPAkbFH/PoJu1eOglFdkD4QKGrFOgY55hOI6av5DPDxhk6DJWDN4
eBdubLPYqG5E/U8igEsQBA2vdB6VWRe+t/lXf0iirMZRvymz9Avz+aumuxob9Z7KXkTKLpgWTNDO
5/sNj3QHipM1II+tOuhTs0yuQGhsEvHyWzgB2DHZV91d7EqqVrFp1482OQoYsP/8QQVZBqhuBlh4
LaXHuvGknk9KZw6IvafVss5JBOIGBc029g9/GlLjOgJ5oFb8EsZnvgJO4JOhfhPArIw85UmRxicU
YV4WZKBL+M/aiOQEdXp+MyaTYiCu08QHtofMLaYykLmNGtezCecCrmTcKu0pAhZXoFMzLY4WtQ2i
TcMUnsz0nOLPCmtnnU3lvo2K0TaC8DzQkuC8b1i+BhleQBtjFH2aHJiCVnOF5Mb73n3387FVyQXT
RIEhUYTL/CNWQ62s2o7BfLkJpbBAqVmK9JWwg/2lRjZeiMLv2SauNLhworjqDulg62rYWXJ+SyO7
2/etk8WGNRztX9GXn18geexh6UE0aRxYWKWEy1OZiyWAV5s2rAc4qT5u7FoWW1Ey1veV71TA4o2H
VTu4LIRmDnmiajAPK0Wyc1TkRqOlUX1PRFFDVEKuCL0kh58UUz1e8ugD2KhX47D/WaxcqwsQwzRJ
O9q/0T5Fd0N4i1awT4xfCxV6Xp882bEaTE82v4Fqe0V1lKf/6BmjvFXsqhUZNDa6PZnZfzmv33zV
LVWeBOJY7g8kWWOrdelQf201NAdU152TbGjzOt3coxq10XduoI/HCsu/9BKEHIlxrUG2twUt7IeR
4aPJvccto3IJ/KKPNQROxk9rNKopjObifnuF5NBRvma3palO9cJtVL3olPtXq8HlvY1ptzww9Bfx
li/VOKN0d2jcQCMWCaJb75JUx8CVO1gZMgT80GzoiUpM5o0VWqKcFZR7F58hQZqxVuNEYFSN2emK
q+khplwK6PuXT0go6f8CQsyT1VPqETjoZT1trZN1f652sY4Gbq6GEm5xFycBpoIuaNeCyCjkfsGI
rudJ98hc4En/3ybgD9Gu0LN7fTHgeWj8SCYROM0QLThyGRxPzGq1kzS2X7Iumw5oVmRXEuUEF7dJ
mr6uoh8U50HQlVI6iclm0ezS5jsJaKLO4pQm80BC3uHOThyo2p510K3B6BWnpNFkr21DeZ3LvwjR
o54533MDkEkLHqcMpgeAgJLbxKl1Era5x1GdBexrScTfxstex2JH1LmMp6lfJufjyAuI7HYUros6
iLlx3DnocUUhV+cg6qKWH18U5ybCJTF0QWxxcOGkMzrhUSmjTKwKqe45V5wOb0HrAGGc6y0TMZrQ
Gh6oj8o69/TDu1TA+X0A5of3HBtUBH737isReATRiQ7Fj6kFSAZnTGCItA5QM3ir0NSqpF4TGyCx
dZlZEnrWKZy9S8mBuuNCD/RkOX274F2IBIcuT0Y9cDdRS1vjv6+wp/h/GCXypDyCHxNGS6qzdeFM
Bm6HTB9W4WbOI39vfMi4ZkLWji4LzyjYDinR6whqbjURs6hEQKz27c2YsdyNIuHFcAMW+PZmqrEA
XtF6QaGXo4unU464lkKtzWkiehPsYY8H8EYBk1Uls4XVS0j+7/ttE7X98uZXd1L/jh5BG7k4nDqL
z6FzrbkbcvcpGTzy7IFdwefvOOGywZ7AnzB8b+aJ+Mfj2Un5x9yoA/FuzJW80tQUVnkPE2IG329A
JLS0ZEj+wtEKb0f0TVCd50r5IY0+SpPZqbnJU3X8YvukpN/4+BG+ymrtD0gKVN9fjfaLwDu2rAFa
QEe2cF3i8Ubg3TyMIyowxEWIW8eRoh3vM3ZmZE86l2u4cNcELVtoX2ckyj4TrjIy0cE2RnOIgKX4
j8uDxhWaTapInpsrFa7o4wk2JkD2C2VNOCm9heGUGE1CiRqHV1gowY3K1478GiYE87w7g4CoC+I4
Hwz25aTOXqdfQPUM6XsPiGlInwbZuUGlSYf7liI7Ul6FVxy/EuOaICkqFedGcBMioXLtwjeSjqYP
nQG/jSkNI0KnxAGEHpGgdzSnET7ufmMCnXTAXug0LkmiCiU1OEKwpsREgL9IpQuS7fDYsXG4atkY
rZl04duEvWA0QCZP3HRL7OKjQj35xbQ8VY/Qr0n3eX9iBGnRm8f2g7AlRQTM/go6DWIX3vL484gS
nFjqAKmy00Y2jch6SQZvoGrCpuekEE9itRhLgzbt75wgg5MPmzDa6DeFuFg4Yj7YtLKQNsaulxtR
y0hy4MsDWH6wCSEonrFnQlcx6SXztoboMWxUDZOsCgY6gK2jeSnlS25587SSMpr5MO1ZFCwWCKPf
hMSlkZj1IHSSNj88IHjYutOwMEJe+OssSxK4cVV8Kt2/EDYeI6c8b/wODsWuc6vY/vnxo9JaGze4
RlGStcoFLgN9c0eu2xoasPoYgp8fe8SgwdSdfHO4geV9ZmFHAf5IxSxuuz/efP3CDrB8wp0QOSbm
EP2v/GkRPYq4/KuzwPTlNg29M06xjY1GpFpHcSAl/suKYecUMdTOzoEmFMaePBWvDNt3UVxm+dgm
8SqSnlK3FGTX2eQ6wnlFyYDkxhknaLKnKTR0NJtwrvEZnTotB+pH6qtbXj7Zr48111h+2fbbKRhC
jHVZDhezl90qgskNcaB15Xt5aAEHFgS+9WPv3H2Q1H/moD2hZysk5LGyGCeUyDe9P1vAELwtXrQu
w313jubx4hWT+IIvwkG3TjAPOelgrbF8KtP1vfVvbKexnTRWTg23WsSbc4nXEPcl2NN8mammJscY
bLbaLr95zk7fSVbUO3fAFUf2kpUnnjEhu3rV9kyca/sjePxnj70teT+cF9NM3fs+dlvsBHAivUUj
HMTgyx5AS1UtZEhBmRxO9U96rnyamjdk5ZEIUhofN7KpDbcR7KUFENVZ+GeJDXohIu6OOEzY+Yh/
7/+AUobCc59+5kVV60NyK8pxzSWP+a2OZjxogQ1wAs1vBiVFIvXykjBlYr/lMkGjeMDvOmitXiMx
EQeyi0mvyh3sbeG4Ux9zU+7Wmk04GXRU8jtKSYxhZAnMA9lubwtVyXHt+NX1ZiDNrvcRgMe/8FoB
/alev3gGBmGXTOHrDwXkAH49uG6WQImKbHuLNKQphYXFh7Tvfm0PfSOz0iYo+zFFQGVh8voMDVyB
k5hn4TRDnkvykmsR7sAtoNhrIAsDubSemnFUbUnPsGqYae7QDRPwz6dfcwFLs6RHA4m8rh+8mFaJ
SbVJaN8scI7ds87jwTsRnf/2+l7Bi02WE1IHH5XKRROA9YcQ6tgvq9GWXsJ36xWKG7IWSwNPhzA1
xi5EheWrDRaNH8aSU793pnzVw9goR08ZTrbF48SxG2rvm7w67MItRfKXZL6ZeDQkXqP1jYV99QP6
BsNvOgv1ee20OGOLgWxBcbQgLpjLiO9fO64E2kyxXGE9TZQomQFlkxtxQfA1TYWdE753CKbS53cQ
gLcKXbozai5xU56RaeEtRMO95U4EdQBlc06atOdk3wYArciM5XXqBtB7VTWrkK4L7+YUP0X9OvIc
av1OVgmdNRA9Va2apgCJwFXxOFaTpgyfewjKUl3Fhxoml6e108+Vt10K2HKcNpyhOZW8cRuwmppd
XNw/uCn8YW/B/5lQajFXW2LaVImHO0wDG6t1zLddXtBzbeYMvEwfmH/ThMANKC35cOWd5IeT71ms
/axTbcPy75dwTw8vz/lU5DvF+eXV4HKF+t90JH5G9HbXor+S0d/0W1uAf/vMOKZjcb0vwZxInIM5
l78lkue33k7efyNnEVfJKUhD977GoAg6I94nLvzpX7f0W93xsK32H/8bJALGTFsi8o33ylfYmBhY
xZlDssTAbaBifCV6txy2dV7njFFfkvA9dNrZyVMpf7t6qKGW6b9B7BnUoPFw5WlZLjFTzkGFqpAj
lBbldIZxoRHPtiOyGm7qtCIs7/pKwrxuLXYnonfOgUEvEoNHofxX1h6EzYLPT9Lw3wwsTANGNiSb
hzLnHFM4sttOiod3sQuL+4FgZgg9h2d2Yk3Hs3wzSaA2ERk85Kq3mgqi1N1PyX+jQWaRv41bb1rJ
LOxa848ocI3u5njg7mPwi3RCnCY8LzBDJduEpbe64JTxNexAiWZfCPR9PXHDRauVOrMId54q/mmP
5GXywKl0+8T/lTYfBx3dNezp03aQ1qMav4q8NjvNfCF3R4shnRENb7FKn2xkf4AF/OVFaewlOuO7
gOFXYUHyHZxrofBCMjb5B/DMMepYgOXcj+s/DiQsov4ixalbezP8R8+7lCpSL2+ciCAT9MvsVhp2
GHdGWd29+xr5XoOfC2qAjDAvG2HKfrEeRdXTyEvSRPV7DXe+GlHIu32yAfIHTElxI5g+T68510tp
7Fcvb3WtjElOntm8DiFzt8ICuW8yLZNWLM6jIH3hL+zv2A5xEikXYp65B2upQVBbZw3yJtpTD9eJ
A6ELfQUcU/CmeXPLZaZ6DNdAiHOMgPXtxuwcxs94FVG9oNn/GoCSpUoOdwFlUkXpPaatPrjlD9hG
RER5ge1D/K1DA8xPTPY4eWtbBi9pIeNcDMKvbBQ5cYyWGT9kXa8EOB70UiTx5yhgnV3Fh05Iyv4/
DJvNq8GPQHdckySkG0Pu64G/XRSz/PY+X3ZTYdBfES052Vv/+Gz6y1qDTvOwENR8PyMpgujBSuaI
10mka/rEObYD0jME1rfDq2pDdF3/lVLZzVUymjr+HkKmK9VW6Mp3N6eVJSs69ikUoPJJlTafoTvw
1TaKDL7/t3/Tp4MHKBgzMdD4Z7poYkzlAVe4+BYOtW8ZVGWW6VvaB6b5BPLRgefLRhX1CWmHFVQj
zXnYzVh3sEUaNEAFJxINrMV9wMyn/Y3HSjmDZLLp2AL1MvsQl1T45gjdKWEzyc2amjKhI/5G725o
t4PvQ5GsI7rMExYKZgLDt3eZei23BC4jQKPV07592mqS4+jGez9/ZT/2JRXM1QyyMZpoHLp12zZD
Fd6nY1hI1xgascS4S88ts0PbBvoaY5U9dP+R7LBKoo/aAW6m/U40lHWVnl7phawieNBGwX8Y3CLg
VMcvA+tPDR8qkeEzzH24pPHwiMsFXktf2urDvwpyiA4WHRhEqdCTVyP6kg6tY3UAlrK0jO+GHrlN
zhF1V46CMAh/On0qsXXMs5ohunb3K8S8vLL8HDq2fpNIFv/917HZyDgRGROXy8iiOTzXB0oGgPzO
lRRtHbdhXR4ebAmyv5jDLYw7x7GFSiwb4rBA6eBYrbNDtBFRvTJMXE+iwMQpQFTW1H2mM4LEbv8y
dc1Ux9JTB8MVA+aaXkGy9WoZzrv/E9YJ4KapMITCHG/swTr9Hdr0ThquaJt65G4B67rEHy+mulHy
GfvxTTO0ECd8RE7gV/VsFe4TqB7xUztIWgxiGCbS29xlvF1JcJfYNJhhsr9gEirmtNxa2iWW3jvA
5cNVKjDAsmr/eO59dPb0Rkf7UvlmZPbLlmrDUnfwGWnvSSyo1YSJlBDzLw8rGvQT5kBbxzMrR8zG
etm83TXO0v3ZYRwMQ7g7/8bmU/UN2D78fesm3dSqpcccFc/LbvExE6o8ZEf+SCJnDKHx3o9oDAyW
IpAoV9QW92N2JiMW5jXX/aezH5eh3CxWQHAs4YcpzTo2BgrDtAfufjVKI4UT+x3K5iMSb36D8GEq
/hNPxs9/5asZgtuClKX861KnYcOGLJ9fOdHMjA4f4Gk15cHVpDlqWj2ufej0OhW0nUC0wLr6BkEP
FjX5/HFh0kQwhyc2qImbrjufUg6PMjoA5OYS53RuXcIoy3rxMlqX0HBjah47WurIK2UlkUtlMA7J
lVETt8khPnb0Gk30rs4Pf/PHcbBmTGpdA0zLTwjH259To0GPO6j4p6n7Z0QEjbGGW4OKKof2p+tv
pLT3QKSRsQm4JJQZ9susZaupr+qatHIeOiunI6RC2+VEJV4e/EaTIJ/ViyXHbvKvLrC6+pqaVKDG
A60dToZeHgZ2A43u9zdSzpTVDsRS/5pr7xUyjHPqqIVVy5kCLkbo2yjTzEIrvhtxWhpZXu6hqSiP
nuhdVsS8l3YPQlerXOOuvTNgjQN+XRLUvWmgSZF9m1cq7JdNdCJnT2FvCcz3iGJ74byh+uL6JfnW
c8wph59C4aJjgHAEwQcgUzZexBpcx2K3M/pNW3cVN9U8nh5HryLu2iyO4XyvXqMDvQKrAEhRqv9b
w++M9AxpkCu/lSwx7ITO1TKWzYRDQna1Z2E8yWvbG9pJW0RghXpmSfdAYSrXLQe6R4vNDo+lL6KV
UAa9ELaA611XZcpJRwC7+aVNUjL4v1uxuBpP6VIlyqQ1HKm6jwCFqKzPoSUBrxOa67QmjNAsebDM
fiNo5UTBk9mzScwlKEbsQAk0h9x69ad8VmJHel4NMkeHB9SMtjVvUp4rUW6mZPv1rElTZeqeNpsN
8wihh+jIQCTrnR4c+GFhoSxe3vDWgfe05CA/7Jq82Jl4RFXZJvtzBuNoB3IkJ0hWE64bP0zxiVQz
CTliUY+tA1RkCL+KZgWq9rSwUSYjUGYj95dWyOEgC+f28hA5RncuM9J/yCvC6H2Sn8qkM1DXgxDX
dYkjCj0wOY4nJd8gK1gBYyhd/JNDtxDoq9yz7o8BTsWIBWSPFOYHL9QxBb7eH2v+sp5UwplKug9/
rjoz2N4Uf1dGVwx1RKXq3VbrUE+Fru6ZQAOWWzQZ9OiRbaw1jtkRL/YaW4HFXB4G+N5XiZb2B5pt
+qwG3cCCQJwdFgoIUs+StudFQhpb/62WyDGZJ14rDJ/5H65fEMvaZSovYZFuF9iNbSLtX8U2ZvNZ
fy6N5UfNA8JOdATZZoc6FvTXtTTzzO0mdqszJkhhglr6CpvqXy+rzRK1I24DTBANQNqgv7dSXC7O
8LNlCfguKZd4/vEngWfRaBvbl2ACIZa9VpyIORZzS+2qxWG+74INyPy5YT6b9vc2u8Ab8f6vkaWu
vqM5/BWgNHtSRwh89TK84l4LkbbwKYDGLJGIIzRStHA9/gCYpMxSqXghajFga4lCOaoLlAe1LVMR
07Wfld7co/utBUrr6h4oBvl+Cj4FElrFMLN5eEmXBcDCxFTGCVB4jA/4Glt5hrZzEDAufjH+6XEe
UnFApj7Pzqpz94CYfrjKrgcZzWAs0WeK7jN0cfFC1KGY6NxE7Hy73RpKpj0jZbAEfRfGjCdvJqhC
lnAH5cQlH7UuCVywQIw24CBBa+Djk2+1NUErVOY3HasonlL6c2MwHD3KE/FxnmrodilxCHDxlNUY
rnPPO59VUGMd0KG4lGwPxOgpGJbsZAME7O9EtGwYMPioXQWIOuLAtZpcvyHmW+PFNsag5ZRn/cNb
eqv4fpOLaWHUVRKQrKPI0wCNQ7Rm47xkf95JNrWWv5uSC94Z/UjEaAheM9gwAgmDSoC/4a1VFF7y
NeawHIlkn48pLG6tEeL3o1GAa46NuQFUJxHqhjehtT+cJXgBOaLzMnfkgH7oX+X/S5ID/fug0WR3
ssGYOfZYVzYGcGSGylxiO4IIv8sN6Tbg2Wyh4R96G+EzUV49I6QRdfED4Gox73QAblLqDd7Tn+8W
x721yNHBjn51eiLcxfHppxljnc0epIOS5NLCjF/H83dXMebjJXq4MDUqgKxkb4495ik4LU6TTSM5
EefEBGA0vRTPlwSgAyV93lCjLUYqBdppkxZja5jURN9zUiWcKlP/vxr4JZ99y/WmrAE1tX6/7mSQ
82YtUZmQpYUo0nCoyuW1OoO4Fd+RSJBIFuFLtEPfqjCSGP9fI4FWut+vnXVk3QzJKZ63eXQ/v51F
W7TzS+wxQiAQowiItmtXqByWIJVjXhMgmDydpXiSMN4jBiB6vLnIKzVSRryMqDoNDRU8EqGbYXBi
V7e47sVnVQDDrEYUb5fR7Xw5raZgiqT8MwHw9DzxQJ5amc0zEFyPJxClSc5++vmTHR861VNJ4IzS
RxHJ8vB1Zha3834gX8mXrMyRxx/ILabhBuLaWjeYnxahihiLyqk1wO7uvQhDzn6xaUlieLRb8guJ
GLnvW+pPIehRPETCjS+nQ3ViaVZ7LKZVmGx34h30gFMhg8dN2B+m1qIY405VMEi6gQMbMeWrZ2ZT
AXYVjpuG9DzkQiIWcJTzoe5Hkmx2VWcBL7wPJV8z68NIKsYiUBKl5813YOr3vLfTM5RW+MLjG9K4
xzOBk98DNyg8xyjQ8TB1gv2klnAWqan2SPeGQnxa646UDghyXdrMAUQiXtipKhhP0CcJiLIIsonJ
vC0HBb+ISkkHJjjQomdmSPrFdz5yeA8/XREFmkj3aAFHSuGhZidXKQz/41q+L65VYbE95donV7j2
muZ/X1YwFc07RQL/UU6uy85pFvXaV5ryVEk/7lLKu46OHNF1MvHQHbp41d1cPn6bTthXaMNzdwZI
xw1nKLBE6gf7bisXxDLnUQBwE9PTs0cfl5kDetDd56KDYmu8GZ3wDJ0TRACt5pjtNRpvh/uSIDOp
ZQ5/N6uCb0jffgDAyiiXA1e83GWmltDVtjuwqYUuG/+o12zp21nIDCPN8XSX/M/OQPUgtHB+w3PZ
edlKPaGBkA+md29ZTeHHXlgPw1lEId9T0fjzpB/JY+omz1vO2Wx1kN1mfKX+iB3EefZqfKj/bmVN
BtYdopWFd3PL+VJFwGZCl2tB2Vw6qZ0y2TvfYqDI/wgWu5xyKdA9u+lzrezkJ8QTZGa5IHqHkmGD
m86CuIXH+I6zDTY8fuBIkC66LQhQh2Bl1W67L0tDnQxBg1I1VFa23cEdlO13iDZWDsWGZsgPBxsW
dRnBpuRU6Q9FLN3Su08OmvIuLCtK7TR/aujLc05dsALUmji3u1t7REu+2PPW6PGkJT+3KArj+LEu
/jXSIFXqD4TGVB0vpLWIEV+5rw5hEhJhxSWGfNlpJV9DZOP8uBa2xPyMuVSe/OsFivZ9znwqr9nJ
+VM43XBViAsxC9z0o4e0X1vAoyUbwH/ioSEYRczUoc4DJin1XHemU0jHEvWjkn4JFnCGRARKHLiL
3QsgwvWh1SvzHwu9tik8sPKictIbLmLVqrZ91MaT9HLA6lr/ZjbnNoafsK3wvsgMn60AWgNt7pCi
9r9amwyPse09meZ88w2AMxtPuI66yZmE6DTD1X9u2T2evdgPtI+g5CcpbbSMqt6GdKkw9BrFnCXi
tjmr3t20HDq98Iv1LHUp5Kwa3j2PuPFzI6mMwHnpz0FCMj056oYavnvDh+b5LWK56uz2vb/ocqKW
opGX0xXG1RusW90V9gPAlvQWey5iHREZ2rY4+8sklvHpBzCP31FKLInLjTMW7Cu0mA5wPyVcX6c6
Z/4L3fLrATmkmwgcfpb5Au2zIZqzcEyDHeYiV/YtjfFtUbYgLDnC5+PEcKIAgRoiLnGpLU6DQ82T
CsDWlA9Io08cS1c+vb8b+vsmTo2dxtjUfVVzBX0pALzoGd7F8XcvkvkkBfS2zRVe3omvlw6wRs4V
B0EMJ3y4sBjexjfXvTThPwxQhPvkyMWgkxIYuDqbbMnMYJJreSyzV2iL86biGAX5i0mlegThwocF
6rDSkpAkkMFOUbJJ9mPXs2LkApITU/30OBPmO9hvEwax4HDUR1Q/OAxG6OO8JcZFWaLuzi94WzdX
rwFzEevSSKAUsd/bb2nidJmcV28ljAdT/PXy33R/5iAHl1o6h98dbx39UUDJV8xIGkg8Zh5Uuezr
0d4iUeTB1sdqANkRSUiNd2bjSpV3WBOx5zg+fl+8Q9SJ53U4Brig1abwKGqJFU4RDFuFO7lldAtC
PRddpjAiaUgSMLo9A9It1uhPqDbo5e5IyA1g5TFAMk2MtDfDVEXOeNmbTP1pLBxYBwbn+SRqFc2j
YQr0oPM1cDVrTaLNK5XWsyNE+Ijqix8t3KK2I9oVTK495DIVwYLKHudp1l5bs6oWzOCdHuDjE5Kn
fXViZj/8MMmGql3oZR46eu6E7zkhYYQruLZxz3bgQVKZVWs8KQNxghTT219qrpsX/RH00rC/UwaV
+hEKwSbjThZYj2F4Xz4iFzMuBXNi34YnkJdTu5KYU5Yp+6gRiqEbxkAzBSzGH0EQlhgXjpCW2Lhe
yXaHo7lsp0FMEfoNF5XOuq5uNi8jYdKe4QCw5x9IDabUUy6ru48rMDpIH9clc1v71UbqcpfH1iwP
uLAuEciFNJ8K88ra0YIXJPcRugfP7jT+ezHQMR+7zZSpU4Q6/dNcxcpcDMaXz9uz8K3j1Ez34bfY
QSQwp5nz0yL14HcrsnBr+FZdIhoC0nL+FQfBoEgdQie7dkMdHEVE1X9Y7PmsrcCMbeHut8ugv7YZ
tYKkSxdDsJN3J0OILuFApOuGPzZmaVc86eoU2kWAsZjsshvVix59DLQhqXoaLXyq2g23UAjzhkL7
uXP6e65Dqb0yGzcMg/bIxtzVZ7SK0hW+jbI0b2VJeuNQfqQ9ogugaAraC9K3Fm7Vk/ZKCBdueQFY
BD/rkLK8U+BuFr7WAwket4ba/nYTHWmC7BzegDVJAorPBPdpMgSq69k7udGrYd60A08EVon+40jD
IImbtjZo0aPRb4wqU+rUxIQcOLN8dyPz5W5tF4FIHWnEBOzgInkytIHFpm+RH4aI5i0zjD/POpcu
e3UR/ro05kx2KPQnl2hNTAcc3npzE8a9N81Y5lNWi4/Uv7AorakSA75G+/GuGj/EVGCH9+tGVaDD
DY4jGHDEXnbpo2sUIVMHzr8ek1JjUV27aIOO2sh+0JP0zNuSJPsBctut6AYbxQ3lRl4mF6Z1yblq
lEQBEH53WnIRC63RhL0g/BhtHbr925mRkXLmfYltIL9+FSjrAhSxqrTiRjCNoy1dd+ExBzLQ1RZM
11qtglM/TBOKKIu2cUVsghWxNbVIRhTWLj1vWpKaDYpaEi4doZn1IZdlSUqfM0KTRa/J4eaBrtIK
wC2LTWyiWc2866a0WcgL1wnySDVqMk/VKpqK+k+5AOa6jVfdUKvyUjru7vyolWJAn64ZNAJY6gB5
IvB4XCQB4W2Is5KVHNJlOAmP4QqLBmApV3CZeRjKxlJERKihOAL15ho6m5DgrSdPFt5RMAPC5BJy
E34MLo8vwyzcmpEoEZc0olmLezHbaBjSPGFN2KVbU3FNUPZ/v6gLJzV7dOkqxXIcBSfGKdcFchZg
zHemd9kQXRBLPBfPqhk087XpMJdD5qcgJnZkozac7Xd0V3boXm+/o9mrQne0xllhSrzUZJXP1k1D
3K6Vo6ZOb8aiOD8arkwC2hm3gX2Qtc1Rkz5cc+qfoe6dKZtdI8ItuGydCi7OFy/Q0WWlzBOTDYjR
pId24/EasWX+KTC6ik8C5g+29HX+6q1GwM3o1tl3MwT6Xw0eZOQzmodaALNx+u+9P7fvIgFrkj3x
knajvA3ScR+dpvQiPkI4fufVQh4aWYyTU+zU75NCwRunomiv5AYTE6WeUsw0MBAMx5QuHMoheOJr
Ijvr8wkrJcAX970orEH5f3njXbZ7x0nIEVVMgGxvQScn3mCps+BXbUtTZLtmPPVEA3ONuTJUZFta
AGnLTqKxbIYlXjtOEb6GLU2U4fDjWe41s2qhgF3z1PX08hkGGG+oTf8UO8J8Ji46Pb05TwDGfrqM
Kpmy8D2reWBdHNXp/NxxqMTOrjA+BVX0F1cY5WwkWxu8agR5w/t+/SoWV5NMDykMXicjamfWEYB6
0gGpnejxItCk4FlKjdw9KWVnqYIDxVELA/evjJM98aafJQhQasKyQdkc5Ma08WF5erUodB8UNhQ+
YCoiH8q+Y+UV/ggKU/xPIhAjwYZh9U7yE9da9R8aWA9MOuiO37vgrn53I6ZCa3mYgQAwsxQlFFyT
BPaAJRzYuWdrT9+FrlPnFAHTzLb3ipTvttPsaUGe9C+DyjWH6jAI0BxDzAxz0K/Qrt99/HHF0Knl
+Q0iK5UbWBnq/G1sppKEnftRk1JqHdowiX7CePKOCPUGt2WJMm1SjWKjSwoSkpZLKyJ3pY9tBZZJ
aGgRtKpacOZZ0Y/niSnCM0ZEuan7i3q4dd/BytDQ+aAOVIOCHJXHCQP6jOSTQO/ofCyGEUUyv0kZ
u1l3TVC47NuhPn92zg8ri+ndCf3R/tPrE8FNLB4ZDB+lY9AQuMJDVFvo6s2xDSSqKFkUk3NCV2in
srVeOeGJJZecP3vKRBp09W8DZ3VLh1v5WOZsfM6fY51fwOtVaJzJTzWuLy9x3CvqqXFeaG6Ur+RF
D9zfTpHAvE5GVKtTBzqfapDXNvPcgwvoMTrbffGwycn9904flBVGJE4+9CDdCAlTYyl5dUr5la5W
4ZUoAG+Ck9aMm8Y0QFKaOgCM9X6sGvv0yY1HzLoANmCRYbPZkDvkf8feMU7D0kO/D7v4zF2Xig8W
1tIxPbkOp7D6tnJ/angWHt0YHPaS6ktpQg1FfO+7KEgSUyP7BpcFRSApVPDlpJ4CL9NoL2lWXf+W
Bz+ljA71uHa+shB7Y5XqP99dg1q13r7x59Kne2eJHo4jlbnUuJ72FRElpNDvuBn6fvHbFCYKydRm
s7nlwXCRDSl8P4ve3CAkrMI+NtjdWROdgiYQAgVpAexvpczqxifXhG6a4gx2RiqnPIt/84xwiJzv
7ghLNPjK6cZebpdVgCIGk1RmBO9gbJBdPgmif0KMn5lzHnMB5Fc40piPcx4FSk8xMMOZI0koGt/x
zdyZ29u6A5XCOOOMIlTeCNygNvSCmO6kDQ8ibuK5MDA3FYB4yJmdb6uHaftlFOhupZZlCOVCB9jj
Cn1z5bI6V0WRl44dSXPb5oeAkkvuspJ8ZjlFTP0PYCsBCvZjVztHokFC+kvCx3mguhxw/4zlFOkQ
f4MeiJ94hkAh1x4IEOAU6oCsMovp7pMG1CYazVNmWoeKBVgAQIc1ExxCsomFO1zJZzwNaQeuU5N/
6M21500kJPu8bN0rPKQnHdm52Fyu39BUw50ZQ1YClMIJYjOK2e3fDvPRFPNRS5cCzt/dMZh4QCRz
UHspIydCsc7swOFPLBcKvfi7lSYWQqZvdZ+PFuQi3K731QW1qWTpd3EIWK+o50bUdM2JamjxICur
652Pn6jsVz6PjTY7mP1UjaPzEGl9gBB6ApJGF6amv+6s4h+voGUNS90KvKZ44wR7sGish/i9WVWM
4+5d2Ge4wdRFD9nVdUfDdKDQzvUfDbOtQoaf5APRa6/CBaqinZSapYY8sgDAVsjYDmQd4fAKhEZk
kGVCP4YQlKlnEcPpAFvHEw/E9chCeqVmfnKspmWTdbjp/eR8X7IsHRTxQqtxVoj2Anuaz5ohYqlU
RLd4a64yNy1SsXIHf4BlpCLiNs88mDO/peg32kj30/StQ0/Ozi/FIXo0+gzt3DvNvC5bJUyopMDc
4tBm5Dq6Yk1ewnie+gkDKe/BOGa/BPvyrxEECDbtWIkbmJ5gnn4cWQ2AVlE2RxrPt+HDStIO2ptF
/lcKjzqAoZUIvsaGx8X3XvjCOxVO9dP17O/eISkrMnrbhg3fBP6c5JMhMABe5E9iWnNNRI1d9BJI
+RI+0IEqxoXQfip+J4qo8h6KNTocQmAkx0vmNOOpqLaj0QMUhR+izIgBSPOwag0a2ZKyzVl2+6Lf
m7GPWIiQP5oKXJyB9aX6uQt5iOzmNv58gm1BT/3jCWb1JGQTxf5H7rNxVNmzPle1HFCJ2gz1BNuK
nZhUHuF8QooZc2JI2s1LAmGSdUhV+OFEkj/kId+FIPvE0oxcF2aH+CpHZAyWqyL3ZIS51pM+rR1p
Lkl7AI/vE433vWUWOjefm5y1T3YJ5ZWz4okV4IieS4SyxdkEn0AEmerMbuYa+d9nkpyEsRd5P13X
S/lNY9bS4ZoKf4omhEynn+dGk6ba7oJh2ht9m6Shc0/qDkMttwZ5W0ICQK9i7oLYCwVhRukDG9Ce
i2taJ6UpxHa/K2k1l8WpSk+MqpYDQlIETV3EBovXoO2uO3PgFMGrN4SJlYlR0cABLsiLYeaC+sh9
J5wareTbxOyaBVffDfF6fT5X+ndIAhkcJN+NRvWIZcqoKHuJOS9mq3Hmn8XhZOwHPIt4s3HDuTLK
Zd1wGNKUaj5GPKAhAVHjVwCjVCsugNd/XCfi5DkjifMonusA7B13KKm7k/pv0NPO4cVu3CVkBMn8
SXo6BfLu8eoLwAGHJyM3FLhK/VtlYwwj9PRmk7NsMQBYTU6DYk5czFnyubQZ6zNVUO3U59G0w0Dd
EYVcNv7oS21TAcctEJTiUvbvfSQw+WDr6n6oMIkGa1eog85f3kQX15k898V5Zziw+4pjE+E2YEHr
pITzw49zkjYtjKsLVnAkc+W6PVib9kLpJ8Inz48tMj93ZfQ9hVCtA73wXNuHf9TcNz46z3cDpYyg
6i9VcVgD9J2y5oP/hartNQ0nuI+wuMBp9b6HkdpAlO8O0zeu59udbLSFU8J75FfGeceKkPyINnh/
HTky/lnMdjXqyER7p3r3lK27HWPB7GwSp0tA0XgQ3dytVmCx1nT8xHxJM9i4cDf45wcKicLot1eH
qvGz+5+SUiDKigQ1MezCf3HQkF8EjAs2n13qSE0nXhbnd/eyEyt70pme/vD/J3irEWWlXMr01Q6P
vvTbJyizljQh4OmtZRTL0EJKHCnJFFqWusMJjYD2Zou8zmf0gvtkusQVpLbBU6FCfiv1jxJKmSOO
2yojjbFhT+XML6tZ7dEawo0EPkJo51NVKDke6kofMsTFqB55S61iI/jEJJHHiqV1/u1uXUMVVEoB
GhbNkmvGMrOE0PAMY7jTrprgm7kXBDk/N7IM3zAFrsL06DQzM6msTit1tx38x0MQKWGhqN9IhRGS
ihir3W0nbbyEsyiLKfJTe+LGhdfZRO96Zfo7lzODz207m0yMdhNlWeMYe7gUwGgdozIx0En8G+pg
Cl6C3ef1g0BQSkaubsR2X5LJNJ1oe/iPcQ9Ykc5FKdEe3V5Dswk1hV/170fMgb2QnAyrufHJDeP9
r+wqt12GDnykpsRNr3QUhfBmXzfw2GJSLoBLqKBuPz/vuq+pvKusQ59gTS7tCwU6cSxs73e3xK9Z
cX4yd3MzYXETzqa9a7uPpxlfhQWQvkGGLYDV7FtGNyhBuuq6GMifTmxyvl5nND9zN3SrlWp7qoZ+
SvU0sDNLZqTkKmzfzoHA+3rGnY33SEV2U8kal5prqjvVrqVuJAgqYXmDd6A8A0m6RHVW+KXINddS
itVunrDx083WzOVcrQzS8qnuDGEw/9JgxRm4ZEZ7LXHW8xw3EO8F9mveWboQfcVCryfRTd+AHZ5M
7YoYkDHRlYn+ZidA+cQsafjy0xy3YsNRZMVcuXk+Z//VBH+nYDdXkVJMeEOBTzjHZDvOBCXE3qO1
0ShIPraZ/ptoWRwatP1Vv+E9Uofx3DtGBIfuNn614ED879VWaQNRUvsgG6si2zxpyVxGAfn7G8qx
skjqcup6z9H7XVTRRrNfn2ScuOPbubmDXEzRFZF9epHLy4WS0nwcZtDUm0/jpZY7h79ZQfEwFfjo
C723JSlkfc+1CicE5cgpq6pxTV4KC9a8uKr2+PIIr5ctlY6VTKLVpQRRVTMi1aW8j02QJfoPKK4j
ONf2Mk0Cc/B0mC8OlTOoR7XW91/Z9XBFLyQ0Dt2xheq5WudEpJOPICGTJ4gud1afTuJkbkFiooiz
DEfaYjgzDlABd0VGWHCxB5JYg8cpxGQVjxlH5pqdcrbWvKk/rvtUWhu3xTeSRThNDtpO+EJXEZvI
eW5Ff+tYn4LFV+Uu/t17cHVxUANN5XXXyYLMafMgoopWqehv6WvU4MokQEoo1ZxtPpq4jWHqrBF0
RnXEF0376mL8vyct3hydKn0GqSjnmAYILGBm0C9CYE58dgA/TiXRUajoREVulIy9kQ9J9P7BB/Jb
NAjE/7MI6Gwgclk4Ge/PQk8dqs9sRcdk//AkXRr1uhf/YIsWcELqNRp8JmKTLiDsJf6MUbbtzw0G
lzT8IhCPSpX5VUmw1HiAqyRI0T1G80632vuzNgCzaiCy2IRYh+Pauiyv6tQXLTI7tvxfUmR8a9c+
o6PZUt6knTJC3NOBovJcMRGd8lYve1t03X+UP41gmnwhSFzRE3pWK4fZZILD5m4ye6NmsSPJPY87
uJKh4IUnpGLj4Y6ty1Y5R23RUXQPJl2zuRMrwVpevrIQ9Wbc7FiKkrh7silFYDP8N34llb5zXna8
IOt3oOtwjaYLbSL/p1ZnOcJNDT3wgZvSL3DjqNkZIdqcciosz245+xd4t0QDQ7d4rUEKNo5eucxy
cmAabhtifyeCHREblvtLM1x93v2wVxIf+7ddNL1kmyOQP+wHyzQGVSjgGYSxG+nKLGTzWIxzp+qR
OF4/KLSS559NB7CcNebf3Gg840fOhio3LhXlloxvzMqaSG/a5ztuiTscJ4s6JYdWy1CXelsUmqYw
/0GXtBs9UgnT9CQXDG2VhzjuaBfm/vAiFyyii5oHcf/3Kp2GNiEF/EZQLzQKe1p0DfIsH+WG+T8G
g/qvJjRdGmTugdm3BSZnbp47HKO4Cyfo83twraq7H9+nZytNVB3I0r6uziJtBllyEeo8t0wNMHZ1
T1mgGcXXxOVJJpDQpu6h5DZS9EzR138lKKqSQkA153t1nKIUyDezy8GagpJs6vaAox7q2cQT9d3D
Wd5XNq1aSHGpgxhbWB5D791PMZsxE4GnjCkPcoPeftiyBh7oYUd4EMptxDQKK/yIjoTRzQ3rAy2j
WDzhvF7xyKfSJEzKddBOO2o191SyISVEnzNBte+HlfEze4o4ZoqEE1iCVSfnfdGxzsuhpEBB4lMc
vtYNGMzYrtK90Rm/XEKaNbtbroMeqNAqXHXgdZ52egOj15HtDoOVBVEgYuoJWhTr3fbGKzwdoqoQ
sU/D3kL0ZElP3qoF9ANXMvamUsql6jK96XkGqzHz+FItWpLT1M6KiF07J7S1XEX8RGSRY4dLBI/3
Ryrvt+FU7S2qKV+xiwcGD6dwocYV8YPVk8Y4Io9z6hqlf1ucnNnuWzn9KqBOxO8LMXySkLxj8TuV
pS9pTHRSXwZId9N0w7IYtTaqUe+9WozPYDXlZaVJLzjw/nJY1NrDxGlAeLEvY8RjJiRpOksFMLLm
5q4eRPsXgqDJHSHo7X2txDvVzm/xZD4nBigS6VQRiVnamT0bkHtxtjaUG/2Ol9rg1DG+1bLp6COw
GqIexC9fJ9T1WvgaU+T/r5nvB//7tekvOOvS2XrW/5QCd0arR2gkf08KLXRoypgWA/6sCBaTpEqs
jwGjpeCjnoZC08nm0eJMAIaFOlVpYsRiUlbKQTElSk7XzRGt5A/9K/CiuaXhpES+fz5TKjka6GNA
ZKL5GtfJsA1x+5ZSFrQ7zvbpjjsvohQjBbUiWqXhvQCwt2csIpTBqZ6pWW+McvkxQseYAhSEZoFh
jviPCMArw1g39Ap6Xu1SS4ZD8xu/faXHREDZHf0TUp11A7qxI26cW5BisteNRwDqWRlRCBsy35sr
nLm1YplfMUFRcKRtDDQIwN46AjKxL7Lk/fSNyLnM9DAuwS/+ACQiQSsr8B06doEFd/OfKP2z+5Kf
ZCUBXnWBTmOyxOlt8iq4uWkbe1BgbP6Q5yWxcMU1I0VZwlv7DqveQCXlaQM0a3+leLI+5Q+NwrBm
XhFeX6xrn+ty3sb8LHiEqh7jYWd4bRlLcFeSSzZa0TEfBSkxbQ9AIsyXkdxZXXqSNfcjED0lnUsW
fif2v6adCfa7yQc8EUz3jpEaxtIFbUPchhOJ6ArBgXZwkjNu4hyhOOCOk4DgX8vzslbZi1/BwzYE
ABxZ8maJEcitXxeDMlYltavOWJBjPv87lFNMQIwyKumqlduiQg+thB7LGD9ln32EInryuggbCUMl
4QWipnUv9uoWsNjBd2wj0Htp8QCI8VzLpV1ACUux/S41EWaU8b+p7gyXeqyp0GQA6mcFtevo5q4B
UlZnvHGoC/JzCCpd9WtcD1PZcyniQLO9/werMDByJzqazJlRHjSdhGSvry6DjZJ+yHcHlTqqzhYy
of9UJ1NVUQsAOeIyQH9O12QyefSJj+qkNkoJSMulzPTlZyBxlqesM652Fdhd3E7Md+fZPug8gQi+
1JH48vK/sFkHZIPgCwbVQvj3y/vEpxsYhKtANrp9pE+0CBQWEcMzPmXnBARAXPM15JYpH1phlZ2K
AyoGPUci7Z3sRE2q82BORqk6bi+auRzkloWeOvEtYpN/3M41FYeHXo9dQnfFl2bSNM94XPNmm+Xk
sWS3FrzQ8dSklLStQ6H3jWzqLXw7imnmQAGQEgGlKX+9Xk23c2J5XmMAW0lPo/1OY/QbNpkGYGeC
HNfO6Svy0/0QusR//QzS0OkDkvQ6l+deCRrb/zBAl0Q5vHjm3RD9ug+grP0tEKrCd+N7bNw4pvoO
FeduZ5DqZU7ZdtJW+35hlKdmXjYBx/r+igiwVtCV4gpcCzQpXhgsRbpPh7yIFST99PnUrpqGN+vv
5nGfcGmjCndIo5tmhzE6HIRUMqpU8rC+jKVbS675fP8l7ParwvmXEe7a2riKVI/+/mi6O0a/h97L
5OueXWDLgVHf5Gr0feM2gVD8iUxspLbIzE1uswrdEnCWuAetmR45EjRLFhR3PJvUGaS9DrHk1qju
caFI+CfgxVxlPK0n75+VYQg3UdFw0TFZj/gvbxMcx2WIy3t/pQhWXZ5oFOZQ0cD6nR0OfS5RZyJN
IkwNVXdxSDU6kbBzAvjm4C568UTsFsgHZZciw37svbpsrKqh3M+y7uCwKhSOUUuKrUqEe12gqTpA
Y0AJ3S514DtZFO0ZRmDc8QXng4Psunfwt3YcOrgU1DXCE+5ZVqeCfM/St0m8609lzW76ZrYjBIdX
e66gFsKOhsx2j8SM7mg+3EyRLPh1sdfCrFQcVMblWKKlLn43VbrpBrOvH0276quSC+R4CiOsf/Gm
s71/b7bcgN2BFOA/dEH3co2Od0koVWX1GNY2FWkpzE33ncpm3uaGqQQN8c8Dtp4mPiuhU78sYoow
W/6XwuZLPhLEVvgL3O5KIiAoR1qGytjc4gZhwkjmQ3fcM+dd1hq2Ej/HleP4SRALhlpNI2XQ5Cd3
KVixHfS7oEWKyzvH5MbjcLatleRrEqu75s7vENqgOErzX6UqaWS36QDdTuvZ/li6R5/QmmOTVkfm
ZOTMuXWczBvbNFbE4pzNZXI3YR2KVfy+EsUH8QHG1sqrJ9JabKM89I/mpF8ui1xdBdhsPUmxZzAe
Ur2hH55UHgxDHSzNNh4iCfXMHfEdRmxm1vWqaFl3M8hwUZXHho5nO/PzXG5h5areR2UVKfUqAGGA
eUmEaB1Ld3rvDdIMKZt6+9VnAlpcPhpFj6XWUDnCWzonwxVX78VuUlmo304cBO26/HdNPU4zbj7C
0nqeHT+V1huo1w1qZkCdSZ+HC019OeJSEM7h4KvOBTgQ+h9yADnKxuATPw57Psyl+N+UJduh8hlh
2l4o9n3SAX41AUzJK1q3oNssFuppHm/ivXCKwuWf6KriXAW2XkROQSlA6XpikaWj0fI/fZHV2u/Q
k2zqmAPGAix+6xSldMa2V4VfgHU8NIeyOrA2kXjWzDYI9pjRzpDKHASwGddZ6oOzd0cQd1dNpSS3
hjSFb+GSev1uwA7n+dXI8kitsMc70vL1xH7SbbtR7v7TMIBh8XZgnNgtzef5On4jcuD4fIlb02MM
JhCb+2Q8J3DdyOUYJ+aUoExScvT0obCtVqdVXGJu9kWsHnMZgsn1O8UVnSUUd5tC7+hIN+kgzU/Q
xNdD/wiskwQN1V8YgbTcZeBJsK1iR3c4giqbezLnSe7bWORjsRYJcS7K6lsrZFcjWi3ug28xU8l4
JnIVQUahQE5ZHOzRgKY37ohhm1gWB1KO4vTWVUpZRHSyLjxJxwXRvJZOrHP7Txo+btgjF8Nn6WMY
ACpkORanHwiJQ2rgNcNZ1Smxcmf5sTxJ8EEra3rKqA8D3C4+2/ms4Z8INlMZPS+dJDVlBDD0/d/Z
vGrOGT0MUbO3+KhdeJNZMGr2850+xR2n15QgUIIQ8s4JDFIYK9j+0ujkg7jF7jzOOJKYbbMRCkR6
3ETNm4pxjpPfBa5x2FD79qSdJtePZTGgOVMUyKbhJnWJBI2QzZNOpaqQvGvyZ8EtflNRptNkHw7X
MNdNzjYJ7IrGXNJTkTQTbcG1qHTIXd5GOujlar/1xMvE656R5ewO3Xf6jv5+KkhqYcxQaSYYQLAT
MoH79IEccjeFck7GXqHzib+3NmsQy8Onte+LQWQGQQYzcBavRS+00a1EVqsh2omfpWSnrK8BVeWY
LCIKR/06IvI7NIcQXv0CexTooSlhh+/U5PWvGwTL8xrdECfU2njUm7D7dIBU9qik5g5XDIPysj/N
hBtv+1Sy1ysQU8FmxN92YZ7RDSZT5M4NDPsTALJeqd3y3M/1f8hJmOLW3kw4O0uZKNEbK8MemLMV
AqUcvzn0bCCfv5T1C6Gc5rni7mqFyMIDTa9C2dwl3pzB16ofyWA0CHjxp5Yb5uYWlKICDN1e+PYl
EI0TDkT22C2PWtK/QlSeLhqXwfNVmjSol/cL2Qp9I75S4QDZEH5XVQ6sGOGEftmyS8TMe2gYhhEc
Zf6LzCIrabf/4yPj19qEAJ6LxfNySh7C41yxHE0NiRRDd+FKjdZNKCMagQmIohd/y2H1PHm12eWW
hnzG33l3Xg6UWna4AUb0izaWfh5ibb2ZipNMkATVoNQeatZq8lTWlfxdkTMZ96NT5Pu35+GpTM2O
vaBjGw6Svd3SxeXUkqzC0IuXat64pc5oojqEcdqaOFmqbS97/vI6zkNfKxGL42VnfTn+fPiQ/rT2
Tyf8tsBtedU7vnwsRaLTRC/kpOnkE5i3W2rxDM1VCmvRfxTmOBwkWaDqxk/sM5rZmDUCJgqtR/Lg
5LafIcNoepzZjCcQRwCygaMK4OFKh79BkknSEWXuDnwzIfcTMBFZB649UZ9/9okQSLRMa5AnHbcY
IWr/lUyvi0Q1n4/jbZWkqCYRTGl1gxXVNG1FZH590uNrJDfQkiWleAeCm3w6an1Sjki2sr7fTlAf
mMHtXQIjDD7LRRsF9IzKvOjQtBdhd4Vo7BF56GnB6hdmoZDXnuwp7tXfLBFBBMTE1AzVLJn+5K6O
Wyn6n882g4vA+AMO22fGo87A9AV7t8ZoorbpdxVbyRxvxzlnGR52VdopzvbeCjumsglARurvT6IB
fUPQpJhQbik9n3lgdYiWT7Mdq01g8hU2f/LQwjubdHCCg+tImDFVAly55AjUBrjzJxlh7hsIoGUi
9vdejLqWO4tPMVvjUs5UQy2EKIMjz6vHJ+zdiKbAm0p9P7sa4epTYuGGhp7iSLF1qtUXlfcwHtet
hLfuy8muGLsNxXYLhk4GZhCjJC7jku4z8jmv8zGSzCLxv6/CNiG9GIhR4t5TMsQcYISRwwWRBSV8
hTXyJ5IvEy7aYQL8fKm1BvxT3G8UlD/aN7xOsmudzAwHTPZFdVB2f1u6hX6VHDlIClG1TcJm2hAG
3/Xq5VeBSHuey/uQDZjTsC33PH34iiMzIruFHCrvz3HmakaV5iUJk5uMfDLoUB2p4L2wAUJqbEEB
ejmAN0dGIb3klC6iMz1Qk82CmOEKbPrBoxvSE5j/hSArP8TLmlQJNxnnqTpzQhDCdVhsXQbYEGhQ
pRDn473LpRTJ9Tw+ZDcOxdyYgE7PeKHjqzu2kB6/Q98EMsUkIraKbHSty5M+UtbTKj0fDFI30JNa
atVqrrERzu4qn4mqGTCroH5nBLeZPjh+fJq3zwSnuH3hYXxOWc/rff8w3C/V3QmzSQlQjySSduEr
p/u6XSwd8zvV/ae2jP6B+rr0bYdOP9v/H7RMI/YZA9ecx4zdE2Avu71DVXAwJTTjsntgAJuowSj6
Cx1WYL+2w1l3VOH/fAtvMeILkJyjWyFauBqPr11PTrf6U4RZ4ESuqdp57gRkZs1aDWm33iChONGl
kHAXM+dJ5JIPOZ+2+HQ2CbT2I4YiFIYYcg1C32nORbM21UaU7tFNDB4Bts0al4EwpO5rdx4keyrM
/AMe7xBOjusqKnN6Mf7u8UhfEhnEynkpJt58bDTT4HXS7bfJAhC4wn0kR4Te8zBfCgCG2wxXiZ2R
Db7dfJ/LB8xAADQUOopQgR9LQzD+ljeMah0AXU8lPcvO8xxDN9lEcArVVXnYDi9vMzHEMHrqS+dx
O8cXlv4DVj2O8r2uJBoWitEDnDwzt40ValL96gyFZVtqfWOLFENrOje7k7jyYpF3TcJxQ1vdMtc2
/9xpbnYq0nV9qcgUxDURu+/6XDO4D7PGBVrFsQH+nd91YkEYa1sSwlOSlbm700ReFhyR56Up3vPP
dnppSLTmbdZFlNyKpCZhJlmvcVTAaAzfGq1+hm0PgqHx+Sqn+eQuOcm8HwTRgmGLD94he0+OabDQ
8liWnV7EEr8bUTM2HSOyZaypuUEMPyJ2mWKDuNRh4QrjkeV6IzwyJHFq6Uk6ayVKfHxfopM7cD48
ISRIyKnPxsLFaDH+2nnCU+QLbIZxSmG/jNG7gXsU+dhC7Lhrwg96DHKXUH1LrTsQya5gRyKseKLI
+m/JXFWcBn6WT2UGfedYnx68c856kGNc8XhcfG12biCJcHAKBKN2SEDuYXD+7Vyd+KUHf0aWhf3G
JBjpMAq4A58VyPkcpU2nhE8UziUCVAi7XT+XlfXWm5soSSjHFcwi/0fJ/vCROVR04XjUEhX5PXi7
WlNJBFxnNc46XugP2HWaGVXY9gYQhHi/n2WniasvYmBG/XWIfuUteW/j6rdzBT6a08SMzRkNyi6e
VcyzliKEcPz9hZ4aCWtxRCbT6zwJ30pw3boGK4LP9/YVgEgXzIrXeXxA96weA2q3YMHgc+3uUnY1
/+0fX43fH7lLEZLW9Wv2dbIsMCy652c3b8UDT1S4SRdUwD5aiDo3uSDmsGFQNi+VZOQiSFgeVRje
T8CUxhNQ/l9w9AxbyOgQBl1FolovW439n3/hIchR6LpBMbdd3rdxLVJa3EXxNvPjkyDZLnLzD8mF
PLT4vEiHEF3j+oCTcpcZ3XeYpLe3OrjWcZ6BRg92V9ExpoTlWxPNrzyqkFp4XlCJU5f0s0INV/Qi
hkMjKE3l0KkcFjxGcbwxnocYhz3iNPvxBZdsoscZtQwC8vw1yXrJJWZgPrkieEfYsJnwIDZTewg3
npN/GYQ86P3EEQjycwztjR+qGN7T3T2lBGQtbDGMcKwiD95pceHsr68HfXQz8GvtFuTbRWQOgVk6
12V63PkClTqY5pPTYwBhMfpgsBL72PytIggW3veIWQaYeHpNynJsDFgDbGPdV98n0WmiD7wQqwBe
IEV66VDo61dfgjmFacTvOGmgV97K7B0melizS8v6sowSbty9U434Y4yT7N+QRx/wUZEZOj1O6YhH
HrDXpapgcqflQcLATGORjJM/z8j9FL0bnqcWZg7gcqhHxN1xdgkq11Rbdc/IodAspnQU5h8PsG73
32c8sV/pYvLcWrJJRAG2iSNOYUlvxaU1c5rhOafT9Nqn6kkQkyB9JqB4L6Y8Bhrb4cBeZAP5+tmK
cNNsVQAMN4UjdnP1tc35kwmdAJJvj4wlDY4SQoykkRKb/erjAjbUf/JKpSY9OSswG+MrbdKPdPKn
mD9sqvDX3BEGOiW1cX8dD/b3U9f8xU65VMSvfP/nwoNk/qgaUPCK8rZ/JN4c7NWr4O8IbSV1U4C8
LN9X4Dlmh/Rl+w8FgjAAI/rE+Z+aGwi2KqOZme6NNov5/6KuG1MC9zlrPVH9SJKPZ/U5NNW0Ixgg
KsdUkLVccJv6YWYs+o4/BhYDjlY8xNcw2m/6pW1OJ6tMQHCMOQ48+fO9OE1UNu18Nd+QQw3iYiq/
GQ0itCGYtVjnBKQtW8bf+pv4VAjnW980sL8RYyGHgTjKHwFxLUFSk5F0wyVfQktN74KRaG6cRkbY
OCQS3SoIbld5laQCbszRnxY3hmUBrjZV8ibx6nb7Gt5dEkgrxJLP5uOO/SO8aMeB26NsXui4aphH
KFls0hJw9X04A06TPjggQHze3IHbNrtSTRl6FmCu++34KX98JoaqY8IyfbXVERxFuVB8zr8j75u8
O3SQV/Wl05aFwaVUDa9H7jrnffxm9hA4DUGZWWLst51V90yRD4b1ZYt2jNebY73laqyrbiHzr7mq
uCIJo9wL+OsmNkt5Gh/pYux3ev6/UnjzR6CXXeUb3dAbGf5ib8UdAOMqnUvsry1TzaZyfJWdybZg
fSsbFriLJBVtNoffHOi9BL1rd+Z+9GA9649B/vvH4TV7PU2imXOnUzCbJwQ2/J947xtjxeYyD3Hy
/Wd67w/kIHjH3DSTOE8iezNqlbpImDq+9d3Gg4EmjKM6oD6OuM2Uxwvil0HLIQxfzjQ5tR16VEaJ
pbUHhFw//QNHkfLLSzjj8mIgHUf5JFQk27Mt3gnuYQzX+Wm8DguvOL9Kq8mlqjHbhm2OOaB2kU1O
BgQgaHIaFURC+5mxKrZzstgWe3oBkgdKCcXcnn2NzMJ4rZvZj7emofTzMNkqfH7yoQf1GxQjT2aH
IJUCSYM5v5sTrL+XNr00utqSFLyv17hV2/eHeACL9O2X6p+3q/6Qk5yW/67ydJ3+POuXG5a9P1Eu
95n3mQoV2qYzhu/QPi6q8ac6FSip1KwoXwUvcUiChSsCkKYWJ1KAnHTscG9nx56ba9MtgTCre/VE
+UDnYvFiH+CLqYCql/joFFffXfU3jGbdXQgSucdl8NFPHlQhYQbm3OWB5i8ordg7bY1V5htkOw6a
iDJtK8Ph9b/U6Ct0ezhIsC5RQU/g/CpVE03DSDPw17sPjIq6DxnY7SNBPPCJx6SlPDXKerSH0qgE
dmrfVk9gWlSYFdG8Sfk5LAPopI3KY33qir1q2cjUzrzhBBIiWcmQ++HhlGVk8+0JfxGCDFkoWn4D
bgzJU8MBE/wHSOd8hPEpakUiNAz/Y4lQuBkmZFud72iPip692ONy/iOnz8SW2dVmXpbxLaAro4QX
Ma7HNwJWcDbW5gk5kz4o82ovr/RjimcbOxmRV8j9A8aA0SmYZiV2HMzSibFbFdXjKai+mjE5p2WD
hJuzxcebt5pDRyoRn+zZXYYCxwC6+myMKF2BB5NUsbmDHi4onrKLeMdEKqJif3sw+AcQhYHYbGGF
oiRkFEcqkyrkSDz94/S3cDD1TGS+44ALBjI1npumG5JSIqxfwMnQ4L6ejgxR0eXFVaEhDlGDHMsN
DpG1D9EJYTVXVupJ2Zhj1f+Ta9XMYqqdjoKnuq4DtfzGvUJ1bb0OmxjZ6zKlyEbecmn14SykFth1
AMXrY+lOufoczgAHryBhAlBjzR3j0MEnFWniX4OWnHoYZoqNQxfJTAyEVavw9rU5XKU05ok89NZ2
z4iOZQSWXRgICMc/dpbgjIT9AffF/Rmy0eCtNY8vnVZN5cAMhwU9XpeQdbYC+eIcf5Y0o8S6KCm9
lwtNl3mGo/e7BJLKDBMnsPBydLtw+Frh+L2HkMyHJw13LJ0HbGVr9ns7EqOO34G32Q/yD5oKXJTU
Ob/+NMY5HHTsbMgYBpwuAOo22iI9WEv9TvOTeVeC3cN0Xp2qtCLMp7O43t/RmPCr2lt9RkRZp587
fMwuQfWAuEbNBfFySRsfnXqlXzteCRMZxFL9LO8cyZJ1wZhxnof5lqRHkH7bvxSt4hdLmGXhAR89
8ojJqn20RohIqBUN2pbopRJydX9Ks2r70LpxEgOSbbWXcL91Zru5MdXkoyu1Y6B2q/vJXdectryx
UKYcElmz8YHhc8RtHKCPZBBGNsrca3w/4580vMWM5bRVQ+5OunEfhth/Co66FIn+Mca4yZv9PtQv
PjEW88C9KWtxO8AMc/m8GzxA5RB4eWQlM6ZPz2m1He/bxkDIhfe/v8herkEQjh+znJKKjgSRXw0g
FT8LSRDtjZioHSX3qetvUzQ5G6BlzctRIw54yGPPzlOLVXgOVbRgSyw2f6t8chaim94NMRDwypei
La0AMCzyfOphdrODJVZJn0TNkFPXO3LmMwRvFqFgPydYar27aNkMHU5MBKv3LVyywDH1A+IzlAhe
bci2tqGZFVkSSrkD87vmH/hHPu1wVq9upQZgMRcC/rkH3lDa7coucC3GxX/qeKL2akxxUOIH8tbA
GoVhEPzHVG+Z7k/mMYMFB4utweMWebaVnvU5K3j9bYFCTu3SEuBo7cf3veG/qGo4UdAtWP3dCV47
UVO5z8yVv8Ek8JUlN4fTiDZhjYpAQKVpH5Q62rOGI31+hFdbMxGtVHOUP6OUQqfrKp8NFUe+9WlG
ZJL5z7FMxOk9A+OlWfyt7ikiuHvfd/k2pE81S+0IfhvPpzneRS4HJ23T1A5OOejCVZRy9If2l8tb
L760jwek45gWAUBqmJQ9DaOQlAoFskS1dlgcuBpvlr5tJidz5IDL3Uc3Hylij5l4YZW4aJ4sAhQ/
huqrKrcPae2l2hhvLfubK7DI3HbfY8w3YS/+dl7o/Dz0LYhAia3TV0EgPEAGIgfZtVqfhiNzZeCu
f8Uuw8Lj65N7pO12dShFrm8kJq9x5TLAj4vfWP2jn30ByVuQrA+wNLvm/IV09GJ1hSR1spe31q+0
0PZrIKGjYPp5b7X7u1Dp/hGHlbjoHl/uDlsmkvJRxVToG7BmkuwCM82Dkwz49hc49Wgy+EZvXhiw
duE3aU77Nm3GAPu1xVTSaGvHhr7mSkQjYr/WF5Mml1u2bIYHS0u+cvOK2Zz3Dn1lEn0hFffi5ema
pYFrmXoNfY4MZU04JJwijFIQJZUDx2COAEeUwNiIFDwpKWnmTpQhYFc4eM1BiexhF2ti/juIuOUY
Rk821KyLttBUip2rHs5Lv1aVO1jUrszwTKqeBOMHQrt6Vr8e+Ox1Xszkg1TT9qSrHanHSj0NXUlr
Ur/07qfKcw6lVQh+IUvaCUIbTlpInCnE6EMdLwFgTS9K2dS9J3Y6zDplhbOGpjcf5Q99zHSRyVgd
vQe7yHfoaBWOevk/rYdCPJ5TIBq7Wx5NfbbEtjHUJy81RdCx/QjU2bNJwamn+gb9gr3hpL1pooJB
wxVo2woCW0Xxv3hMC0ZdyYHAA/VgyEOWAHDYJpld5aKcPYyeNNa20+O+dmJindvQLbB+TswaPwaB
N+6J8aCxf9pmNCirYbKuH+7+cDqJA5jC5Vq6iQhuzNlKIWKgddfTDh9KHDwXO4LCZYpWdtmehpbQ
42iNHkbmeFiwzXcHdRK4VZ8ExAHZZGdenaxTTPBKuWbrr9qSHY6ztXe9Fr/hxb7ZHLeXT39kqmgb
dWacOBzBAxk5ipdSQdbH5U82minunrDOaA/F10I0yv8JOy2V5z2JBGACz/DiuKBeAZRmgYIODDfa
nJ3ADB2oyf4yEf7yKs1X1aOdSTPvnxSC8PW5P3lPrd6yPcapb64No0ek4dIVH1iXLnksWU5dCyOo
lZsxcguOy77PfU+eQxdQoGZzYpT79kj0qFvpDWkdyugSuSDpUK0yTPuiHCzqLNngCZsetUd5lfzL
NXXMI6AGh+WDyEXtDuDvycV8QT8VqdHWpQ27F0ZJshOAw4nNZgr0TdJJQLD7BYb4l5Nu23C/g6t9
7guDNnhL575dCzCab3jAWPDqkRmbb8sgHba4JnLwWsXMq8Sxppk2fBhT309QfOey6XUvQYqNJJZm
3NlIJXbpcsF59OgiG+kJssncUniRZ43ushe0XgXPu8RbHr6vjJxqDld7CU9ljEtUHkFTs4ZYCVbW
wuKwpQAEZ6pURZt6Hi6GqaQ5LdU/Z+28NR6ZuE6hm7kK+XbyGyqGxV+MhxmFIjpGzxF2G6zVAAzC
IaAaMsWzZ5g36gJKp09YSpYXawCunEdFBxcJfptuClcfpPNq8nuGUVdKItwDwzNo3HA5ic6W0qpM
PxEHpRvbTsXoxs3IOO09cwrlD1S9wZTDt3fGkMbQqfr3SId/BVVvp1CstMj5X01l62SX5+s6zhjX
pBUD0UQDPHdcObRko43/8lrkLgoQgpGxXwxUP9xwoJNGnk05odmTEuHn2hQEUw0c/c9EtcQT+rsO
NQ9a4fLHkt9DCRVL9kgyB5Wys3PIHWp2pco6HgPqov0+ClCa1AT0VfAmyhh9yE2HkKQ5qquaF5lQ
IqqDgLNb2/gutvUKIsosnLoWydqPIDxqvb1rCC1H1m5q+5naLdsykcOv5YqDjDfN5U5GGroRUkQh
jOT85Z8AAfXPxIYGqdYj+PpWSa7KvRcs3mxSkdoK8ISksiHv/BAMqOtK5kcSza2qpn5HFb5BlIwJ
cGz+FK3S2S+y8QtC32xFOrByIXp0DJ7szC+2p59lHJCFhHMV307u6Y50uBoHiEqLiIg1lYqc0fZy
L5Z8Qjww+zG9un0f7v+Em47exbp2GC7IzPBAQ5YmyTjzCKBXxuhm/28TFBpwM2KwdGTrQc3VDv0h
SGAWDUnSUybXIDcFevxJ8epbgvdUgTXJ3Yjtx8dCs7+mkLiuOccqL+Yjt3Xk/sh4zQoOcwW/Q1wD
KvZs+iAJQ2gyp7DudtT583t06Gacdu5a7vtbq9QTjhfBhGhUzzu1diYDfSejK8BuC56zWq0Ws0zm
p8z5RAL8ce6Z+PRgmRnzgZ/xudErNOr6q4qNyggDK5VtLpXam4kyGdwf77a82YGxHRd3SOfMuh3n
56LrJH/65rVAl2a2n3jifbbKpKnhKJJsE8qST3OiryDSt7kmTJyyNtMQmSAZXOmefxzNCwX+u48D
14mDJ6v95YgEnDUcBwx1ISzg9hcNkIN4g59AYwJd358csUKA1qCwyy7lCKhWHxbli73Q3CzzYKe4
2mrmae7kCxIDz8QCVo/6AnPtS0tJSJt6HLdCigaQjXONQ85oiBUFT7psgzeIXpRj/hUlJU1dU/cC
wHX+nJB+gwg7b++SslKV83f5Bci0tVDmZ2ccw1w2/t2JIKSTAF/58Yqm0TG1QAeAcFZ/XKr8tFOM
/Qo5HvGXagHQU9qo0bYtqILuOvy4fBDO6pPhO5srDrmz+QaXEzx4/VEUgmOVtIgfzhrnSbWLbvfV
NDCDP16sMHffL4dUaCQvGHmgOO4fmRQDcTJhaylqePS0rb7uW2sB7I/mAhc7sEqeQmRHD4k+DqtT
g3dtBsWRd/5QBSUkZzQ2y25luIBYmivpggdrQRi/rOIq+Sk+tfMo+zbPrsY6HM2c3PsFmhHdzwrK
ju7BYC0b7xBFFicAF8BpggaFA3p2C1qkJaVGAZZAy6BmM5DTAXnKx48fNrbcPZaIi2dbAGuzFl+h
VMlmNl+0gPM28goJsMwKhdyAa0koQmUaQVpiF9Zhx/MCgnPbI5JcSkJQCYQa4YENfUvCLmNL+j1d
jg9nbJa6l/CuzZ2CChVnG1ZwC6Ef+Ws9R3T2YgRsUOaEArFqkoi3mYQqF2BjzEhrJ2RVWRbHbzDR
dcP2gwnWLco4UtPMxALNdUJrXhho4bu61SVjJx71Ft5MFt6kmf/9jCrDHFPTZugOtEQOM3qi0e+a
SFrrKVaGzVr6doVNWD8OD6siQyJNOzIvq1P+uhVNUocfsjL+3iK9zAUGSQLjZji8DD0vdJoBJ3Oh
hZkXvNRc5v5a/H29hK4gh+yslF+2eqU4K79ILHyIci3eBXKLZgz3EMbwX8QQNtcQmLLxLCXuh4qY
FOVUx2FJxb9GBH4D9cDevRhWEAv/znPYEZUpu1D9Vw8U9L2Tvaaj2vndfpLv3q/tMXhLI38yhnSI
XlUb9pMFe1Eh2ZqdxzPSgQ+/7+hI7itxFAdsxDzc8WC0HyydVBYFKGxBRPrusR/2/e0xMqpmJjo5
pDT/fQyhGO1pHRiD44TrkpS0P8W9qWLW8ko5PmMTkNtlpEgHznsBR30b4lVBi0kWY6ZqaAbif1Lv
oebhQFVQ/bvx7mJDOvbv0RGP2ovpp8xrxNDaWr80udBDJkcSDGHfk3VwRnpigwWNTcAzegiL+4kO
/JDt7oLHEK6PFH3EGneQf+mGgbMLmtLsmDx95ZPAVPobH00S8RkoUN78G/9FAtACYXw0KP3wzNKm
jZTmkPQDCwqcN198JjUCslcDbaS/0/MX8GDiEQxUy+syYo8bkvOUDHXxsblu71AGD/BKqIoVFCnz
LeTaJ7w8DlrQmJNiQYIfZM7M6HKdWyr4jerCTFWAE6RNmSYPp0rSUYsf/mcNew/XarayBNpEabes
od6VkenbLdotJ3JvPTAqtqXAz/w8MD/fmxCUiSsRU1qelxI6JacuV8LybUlL2hwVy3gFPSFapt8x
ZzG3+rDLoRqDMyl4AwSO9OZBvfq0h63RrkRC9YtSB2PZMyuBi0y0ZMa9vZTYzHMVeJl67onvO6Km
CDg4WDeTL53YiHkgUhNDVQffZD2qNvdP3oabWp/9zyjAbItmIv6wIjUo3fox33Y3hXbGcsBRqXe3
1HpwU7Q2YExDXb3fScvfETrnFJr6QJR6MWKAjNHNmrM5cIT9RMl1iCrNev9sFZb8hrWgdJmtHosL
X2FGnAcRapwWD0MSNavkEMi1d5C7VdY+aeiqk9PDgGlhHUar7BIujate7PESR8vmMo+NWqqUdJPY
hZEFsh4J1FhX3icU8iR8fXqR7zRskWKvQ9ho0+wLBWBKPJUWJpQFGu4dPQpY3ISlSqDoJQ3VBWd6
p1hz/AcpRV9mfwoJSsogCzD0XMGA4dJ9Tnn4PpHfuFputr9ApOSuE6EL021siePhiSHLJQdkADUE
x+vc8SSRF93nNMFFeiUC9gZhelZJpXxeZxjSfi5+o+4S37Wgwatan0OrIFmXKTTbnLyWjuycKSIT
OT9juCHMb6js0yIXMNKCpRIGPg9O6ajuxmGgCT7g8/7lE5iZENoEHpSbzbtPUZgPh2Ut85F6VclT
CozeSX5J144DO+wMwbSDPkT0rDa9MsFw1log3ADF0+uopDjsjBTMAIo+6+C3IfzDT/7r+MAKAADh
k+89akxqsZVzw9HB9vYg0iftzP5ddpShNmm8oqtA4shtt8/LvfKCP4fVEJJjpHpzHN5e76Ie829h
U3WiDp7ZYg9LSVTG/XgI1zkCbKVVcJfZEfHMyQNtqkprAUVroMkaZG7W2q/FH8A4jJM09Lj31QHA
LyScJ7DmZ9qbDmt8Msk2eRffMjZdblMX+MLi4Q3NRWGHST89mknry4dAcu8ERo1KpX8RmtUZaF6h
CUYNo2DFQ57tk990yRn1oUOjDb/8wYLgfwWv4zY5ku5Xm0lXMkMcMNfFQVffSg3qNluh4SjwYAj6
1Thq21IfMgARsiWEg2Gi4qT+gCGbrlBBUWTh1hIKqMc6Hk10SN8eUVmaAoFDopCYr5i2Z/reUu2C
a91vMYDdnruBzbJ0xgJ1Qt7WSDcYLUDLQc8rsOLVpwQ+KdLi4nBIQJ2LvdAjWRksaW4BLdag4bCC
1mE5/BJFbnFLicPJIgU1meE+9w3iNFOPqOTl4HTkwzphdsL6P8NbjXjDrmAHMChJ3WGNaHefXc5A
BqXxj6FQVckA7ndqlSA1je37MT6UAcJzOZY5UdGj/PYsLrz1VTs8A5ICezcWxKvlvULzTy58PQg+
ln2vMVUJv5xRWfgEH2b1nE1tGLnXj5OMHSuXCk8o/F9eEzyeUsh6fyA1YAgIarx3Ts+eOIx4UQ9/
izrgG3VX/Sh017cNdehmTgwyVthR6z2sm2o6sajzkJ29qAtUaPeBH03YwrZPoo/doxDw48XRVKKn
SboWmyZuxGTXBLQRnIXMVyheTO/nw5h5YWHhpB9pXjBuagIzZaSvMnmq+BrOmbSuzdVpNOFg2NrV
I2d/5ivnt2QWJgmLxF4IpWPhxeZTZiY3KhFAeUVS0qD4m9CijPELuIlJA0GuXsMqyMhYjIJrQgMc
VYIaW+pgVHhKOnU6YHkaQYo4psuvfj6vSFXAYGh0+FN/yz+7V4gU0t82yJgt28VbhLoISuUa5FEN
SL9bQVEeLP1eT4jU7SQUzdlyySAIwDI3iKsNTeKQKbqML7xOMWuVUtN+ZKcM8G7EQ+VueX1xYuSQ
p+OEkNeCS1lcxy6njtM0CZBmpHy6pqu5ghuAwYG95WajisWNFf+XpF46uVLWAuxz+U+2FwFgWJF8
ZQlOZHYBpp+2H/pnXTmgK3woYZRsLLe73Y/XO2XARC2KpOsJtx3T8VWGeilmzWF2ZqzUJ8lC1IQH
zVDgCORthKTbZN2OtlVTLFmNGv6py+ZXgBE1+BCiWDuI22fjDNfFTYJcZpc20WJOnVgCVf9xYToH
PSfR5Mo6RGYj3had3TMxUPLFcbjxn4VTTBNrf+l/YuM52TjYlq8osoakxUaf8olQpBEZ711wu3us
ftrwijB0iQyr1IrxF/5u97zz/Zhgs5HmgBaMS/AkhVyvoBAR3BLVy6XHemgEEPdnLLV6uBtfCR7j
zBjH9xFyeDjja5WgaX83QXxcP3tGeYNRHG2z9XEgfKLMU6KNr+d8wKFjii3rJux01vVvQAapgUZ4
OP50eZoOHBmrRggeKi5lxPmedmVM9aCwwHfrdsR4uDJuzZ0KQqEZNWLYT1ZzjtUv8BK54Vg6iqzk
aOeWya9ipwYgEG//KIW+/P++usaZJE1IpuGxNkVU3oj8biBwdzr1aIxh7lCwtgNQbQ14Gv3uJnSi
RVnR9dL7pptjw6wSiftoETnVx3NQ1T+1gwZ++BdJTAUl4sz7bJ1ql9/eNDinPPInoLQWccw5xzgy
u+cI4KqmLY2PFpG73k94pJk4P1bY7zCEY4brkyGHlOmqx2uMOIUGMBKZmUM+FC5vs1W5YMDNBcfy
b7EQgT24DV67BMl7gbe36DJVJST8oUp8qFMb7Evu/6jfm+hOY1WqjKQXD6tSbVDPZVazB1JhG9LW
Iis06e/Njl8GIYlXvtIyI2l32Owk098LQyabsvaLlG/LqB77glMG1ojkyVgjh3O+rL7clSoaVv5M
qNnlK8JXqe/ll43kmE7I5zhl/S2rOdspAD0zQAd9p3osM6NXkAz7D+AdLtrWdeoGGd0oSiltb39u
DpPOWPRu3thWxTdh1SRAU5ah9PAS8VbRaY23ovVl2e8QDtGU7/DdzYWm6cGQWLJnk6HqI8BKvaN3
itHSEM5BySFTF3xSNc4NlH5OUaAQJ02Ezcwin3DdebklYuHMg5z+64ZL1N8WD4FZHM6UHX/Sohys
LrXI0B813TLABkHgVAb8YWfEMjtusNVfBryItZtdY+lIocm3ljd9KjHppphTc+ZIcgSnicmEjhJD
YkxFvJssJ7ckAtCLKGLSk4qBpyR1M9q8IgQzSl1JYRGkmoNIN0Ftb92wLyXWXJiMsBs7bPgXwt8E
F3il7QsjvdLIqHz+4/wsyTM/V6oJN3paRP1qk8rcNwk0A3vfVGp3yQbinqzVfMG60l+x3zTSS5uO
BiMeC/G7fh6UGsSceuTaMWOLfXayGObYHKZk4JDiPYS8qU+6tUg57+dZ/jI6ewwaerTcyKAg9/7Z
tnVCUlBqvlpRJcPKeI5wkcheoBBPgWMSMGoTCBgDnyZ7xkUcSwLZTwbu7sxomqzNA3aHmHnhpGoJ
UfimGsGLrtIYZdLEbpGGHwbiRTvWCAHdhTbToL9pR0jH//zj0FUcDKDKty/hmQws6e4esd7cDMYW
gXgWde9Us/QUH242+0ETT8XxOGdxfibtGjg1wdKYc1diKw9gw0dFqE9wHC7rII1EsgXkhyfSlCFe
u65nCYNw0DZL17PpQrIkpaJqe3/oX+hvnzO+mQbs1brF1ED0BmnA7VJM+uSv3SkMTLfFc+itE4uJ
mCJSp4aAnVDISi9JVa1ql9W/NSBSqcNgnpcaKQ3vUe9mDSmAnHCKBrVBDRtQ1vY5MDxXSrP/3HOG
qOZyj+4l4quxynNTNpDiXhe9/mrCURFAu7ehT++mTz4ZeumNnNm76r/SpkYCTTDz9B9ud2WgJF5E
zXd2JQ6oLDxkh4cz76ys+ky1M14o1lhXkFdsJqyov8d2idgDNPVm9Bk6fFaKH3h1d0ZWbLihylUy
XX5EEwqI6PVOwv549x1dWlvc9439gqpGdb22jK4i3JtuPQeP6U16a2qVDJWVVUtzDQvUTr1+Ohlv
by063/VVG57utN9AYtfwHaGtTVwsVgGpSraj7jj6TQ+w3mXyGgBNYwJCMWdJ17eAjX4wTAjY1RZG
hd6nLtnlrrN/lrnJLH19NBppTqMYFquCm4gwaKydOOB77ndN9VQ1mXyezjMG/XTRDgcAJrNhl4lt
s8KP7scgcTiw4un912Vp2y3vTvy+ME5OpS6CaNlTQwMQj/XPXqxl6B9atsL3DoR29d6HuqLTaoGC
7DXD9UazuPvEMyJfd7HaNjTl1aeacya5+3jSv2kNrj99qrZP0P5A457bnSdtFTWE9QLqF9LZbLyX
PtSenQOf6ra0/dM3mGVFr4TXLC4hfsg53UU+fa9K903+1uyGcpn2WvlXb6QI5Qx29+Saqz9Vb4YB
oJ4gc7boW2ue2JRuq1VMjS2odcIDlrhJ0cNw8LY7mvlAeWVrXlLts9Y8PcctecCqf7Naa5OLfms/
C5l96PGVsGMR0u/mIJMdlOZJblFLt2ECcdNJM22clWfOoVGF9A1Ya8PDmJkHzy5ZOzXFswK4IGTD
Q/peEUSEjbrkSl3MkQ0EUuoMkZUcTvgZJtXRcInUPHC1p1f52J+JqaquqY6VPDARToxOwppfcwqp
HTcqjlwkrCYwFs4yBpuZlzhACNDmtHN4UwdSy+TviU3RNEc0d8DOQvWXIM0q/gyKcqfCd2DNXdlS
ulwl8Bwd+2ZlNYjFWelZuDfhVC1oo5uvykGTCZwS06CT9W11rZwBzVqf2dZWkTEa3xg3nkTb3sKE
YvrFqlj0hhu2fkLhP3dgTyPNf5hD8vRbjdnol74b/Ut3Vx0u/C6W3QxDZcqN6q/4LMj/m49rbojt
kMGOtV6pLIqLZGhkFBX/RDFNo3J+YouPQ/KapZPT9chyYT0xlGCWs9Jjy2tOK/e69nlyhQx84rlV
8cLkBIz0UbpJQJY/HAR/k26+COseaKYMq3toMFQb+lT/yoyBG2Es6Jxq9PI4bHBMiM/j4CvuzPyI
68+aPlLznNpvqMW+pKH7G7PtZbu+lp/ZhppmSIBIG0YCRbw+Cb8tTnEWS2riGy4OEwKvIXbx8gqe
Y5b3Ju4WHw7HV4RgyZcBCME9rXsGoQOo8StZMiktPZs49mfkmjwiHzM6Nm3iLrLs1mnUPTE19sid
Tg0AASuV6bviQx34VQP89WEp/pUv5cXxKls+Igxteg7TP7cvwdIFb5Ri5mOOK7gUQBz1FsKe6Qcr
Ot9R/F9oSWXi7q8jNm2zcOxF8DCWHAynVYxzMMzHI5G2qCjccbiN9LOExvVAEMghv71MBTH+JLZS
FgNXaU4ns3jN5vvyltvrwe+g4uqdL2qqj9JfpPumVeotJiVmp8Nc+PhOXh1vpCVRh8W+3J+dK4HI
HNTKgzvOM3nnBA90FQaPL3KzWLZg+D0B+mSqi8a4R27Q+7kLJPVaqRksJkvDSaetEKUeVv5HdCII
Gwi/+88Bqbxo+O8nVvEQLAz3D7DiWr+VTJkcdqbzBrXNXdPL5VoJjWVa5Bl0ujB0V/AEP6udgFxw
B78Kv5xOZBjgcwrnITNsEV5PebvWkZ2qiwztKWHC+isI4yQnrvv+hzHEXLMVt2vERzyToVfg1B2O
hstlRjwpZ7fIm3XFPBvuY3xEtv+qRrXNvsefxFX9Xh6OB7lPYTpNH9PNuz/9LJlTQFq4gjb18KTI
dkXxDZKKiyVDJH7x57u0ZuTXGuDeDI853bn69u4F+Cjms/EYJQMwKlei+6SnUHh1IVyEUnNmQp0q
TgY8l3E5evdl5mxQ7o1DLyR2R6WnEDnS/POEePplvNdmm2a1Wgy7ZWwHtuvE44a6oF0+p+GDxTwz
BUa9iU45AY6QEUlRpcfx9CfGrFtr05nyVURSpkyixef1N/xWZEK8v0EUjQkMqCKCRC3QBubfcods
7McWSjPkcIs6OddwMHULB3puLAyZtOdRYVyHFPXyhoOU3Nvf4ohIbh0zURioDG3uk67uUkNYTA9O
JlQlBmPAToiyhQqYOlmkMzIaxLv0ERjRs/1N23JWkC2fSw34cQpHqYuNCe5U6E+XkWYm3JHgudZg
MRRqKfDFpggylL/W6eJVoF4vMCS2RuF6b6eU6NBmHwmkFqrR9Lw+/sOW27p+LctUNgy9BpH1rV9Z
ANXUe0X6ixZRsVNWRjRe+fa1SGsjJb/ddtYEfZX5yrT84sr99C2ibpIBc3ykvFJblvwpSDMNd5E0
V521xujo2ya5GItqnX3KOdsAgFSfJircYaYts+UsgHpiL3DSe+FPQNBMnGMq83/ZP87MqU5dczGP
UC+ePlkPQEI0n6uOZRFY21tKH6HTjwVoMKb+aRQQ8HrgBVBzayBOBKbIuWI9QJw51e2YOUrk+bwm
0wK+h9G0eWVY6vf1MwplwUGvEC9wB1H3SoAAM0m702NE5Oee0gZ1hvH6X/oWpPcmBaHc4Gz9reOq
+9EJKxq+HQC/dDrEM/rHZ9nQrivcQwU4OjP5nKAdWgBPptrMn1euvE3Pg0G2mVJNMFOO21UhWz3O
QDgm6jgHptHXKSCY7sJembU9ZdRhFqr+iA2mu01hIQp/P7ZnEgGWQA3d+AdlmrZph2i693Pz2Oem
nTK62Ic8iBG1CHcdAuOYH3+iV2KQbFxJyO/zrAoG3viYx2w9hOuPcrLjcmxpYbJmBmIUWY71ceZ8
wvSyIJUnb4fxifJM1Hwtm1ljgmhEytzoQad1veaRZJqtw2DfeCfgPUI7w3tj1ayLyQ7C77jZdhuG
Qn7l5OUTmCTL1j2xoXYiQmQ0vlYenWRImpSmhkJ3WcQonmLPSatz3fIlES5e9veH/9n4QfcfBxT9
z/86XQ7HJvwAitlay6e9/df5YZzwu0v0wHsBf2XwvSuyfPfk2ZjnNfOwpqHPLUjp99BikXBpPE1R
Ndwta7qAZgOEHt7VIJ8P35vQRwnIBK8AWpMV9tPjFSECk9KTuJG5KqoFWOQVv/Nel8fsKJHssusn
y16A02/Mc0usVZ7hAVD9vYlOMz+cFDD55bYHzLOej7JJ1e80fyEzmVMjgrz3tK/BK2htHWKxsvdu
fHzDISz3QMm4OLg0AuNyC9lD1u3FzNvSyrpDVi4Dxe1S14ZPMaAeaszH86HU6/i3Sftu3dv8S3JZ
u9GoJV6qzjQGx0mI6/xoe2+dMvB4ExX6F/ejz9rucxBJz8E2CdFCYT6Yc9/3FlL1KGk8VmSxw4WM
J7keNGZpBlnuuTw9llzvM4qa320joEPlt/yBqLKqOJCPFTHwSq7ecd+zOP+qEqjFAq1PSrX2Ayub
8cvJSZjMIrXn0ovR4i9wak2DOnyljCtdEMcxB80uXhWeqQmbK5oBjid9nl/eGeAA0DNzE0dc/wtA
4IajRw4UGAIr26fUcE/OlNq8Zz+t7T23K34LffAIjBgoaLq5GobMp3DkW5Ld53Ohl36OX+F77kxH
DCywmejp5vED1eSpqo2+BWOz6RF2N94Ey80aleZmdlXdBZ0z1zM7/UUNAFpldXp8Es2n1A6iMs9S
4/HOQWKDcqynYscN3N9ci2VW0W/+wCpJFpDw+Tufn5tWRYXrRZx/eP7MQJxY+BFNaIJQGYoXA9Tj
qNhowElhphavWKew7BTmh1CHTrgU3geGFuv/VAqeREqmRcWQS8T44gX3hvDd3I23xMBxm4a+AEvO
7ezQxnKST6FdMsWgsnNj1rT5flaNZxA9Yr8v2TeRmH/6Mvw8vK3ZtHyEMsI5REUolHqsNUz51NTN
H13cTqWSuLRm+9u29HohyTv7HHw5f5tlKgkLcbxBosgcF+O+JwmiLk/DmYN64MXk53ZcyEO5LjTh
cOQbs/ewUPQt9qBNwPnZErRXbPY4vSV1GcnObcZMrpB7H2L7YH8gPCpSeG2u+8g9AQcJ85PVgpDN
YGx4WBIwLJfUQBf5y0KlaJYHopWz079p81V7P2onqLQL7ZIvtYOsqOslUlrKEyGYUmENO41rRwcq
siV+LVHyQNbRVW3Yp6bZpRvXZhklbNPwJQov3fwg5FJ7zVlP3nnUF9sRRUlrXQNo2rm6UW8ulrIR
fHrEL9xyIwMylYokWwQ+cLmng+MxKFpDm+5PN/EyZRe9YfCJHw16n3tu9UtfwNhgzIFhZDoVYLuI
IXA+oTM9SzAA1nJaDv1t9U9wEJ81FArwY0pgZGit2CR6NMKJCopCGjPjAN3uFGemgIetCLkwUWZD
JMea9P4KOyyQAZaE04Afyvlsm8rYzHKbDanUb//RKIyXYpQlzyCyQhN0EZaAymsdC/Cy5wXMRqvR
ADLwxPdnaSvtvR4h2ldPjounbMzqzuJpEp+bDozr3s5fRAQflYEAvwFMnWwKW1dpb08dannZIh4e
viZXAldxazDl3N1PqmPuKkW6pq40tt1FQOQ6wGabXanG19c6VNvynd7XBkTDN5ulqNNm/nWZWizc
/m+gBnBzSp1BhUfQyz7EmGqaelv5t+kwc2hj0D0h7Rr36wqXnDGe8oTjTND945uewE6tMw/afmQH
PpAvbn/7rwX1yceYZyy4D0ATz6LA5I9dUGdtkLN5Wtv3TFSsAJwsp1B5j1ulIF22e0vcEmQGt4hN
wZgPku8yGCw6qs5ud9pO5tZHJNGTuH4QsxhARO6RRQmX+GKDPPB11nvUV8/IxH41OEwKhTJTYEZc
qqlp3TbdW3GSraxgl6b+6ZyyNxX76s755jiq0enG3c3fLUOZesq61UjQfvxQ6NEKuvMMG2lX3jGH
qim73JjWqABd87MVLMZXMY4kQ9xn6yaoFNQNMLsv9vOiOn6aJNGwe9EAuzYdMEnLCMumTuIx/2ci
HFcZt3rdB86ll63YyJsgZfKHF+LoiycprnWeO4i5PysT6xGBQD7pBJ4c5ZkvyIdGCjrqxpwU9oYb
y1ezqiN2dS7FW0B1P9if2oC0LhEBxmELfdnM6s+OSs7TPLI1bBNxXT7gRJB94g/+ICft5/A8h5Vy
gPZ6q2uif28Xs13PeUp2Mditly5Vg37B2+4/bEK7vchmT34Iir9kMJTwOEpxd2UK2wQllclf8h6n
pdQbP9Sq0hXD007jt4FhkWy8opS6ehwmLz1ZpseCB46krlAC6hTGDEQR81lzu0R7BZ4F+/ULE0fN
e8ROPq3+wTZPb9NE38Xx1PpNtNdt+Ppl4fUMmnl8sMhpHkTm4Adt0gyGvSnO6Eotxmu568f64p7x
Kj84U7WywwrSiGpUk25J3ab7m+WXR5YRe/xSXIK8+RRcagRMkZxAYjPaWwIIiw+elXQ/nsPtjKJP
SNjPhVR3CtB6CkNv3rKgNSt4nK0mhup663apdBwiRGaoNr4rZIhwrlOkNSa8HySFmg5yLXk47bvE
hjlVL6+dHA9qGLaiQHw0wtYJg0qTrZBX7QAJ7iZWPVaV4KAN2gG/EqBnos5QKtFr0zUL23Fdwh0i
HXGPYmwZ+/iT0zNvJLYl/XZZHNH/6Z5tJq/1TsUArHbVczn3j6hL7uRQVdDSPnFg4x0VSswdGIvH
3+52qvsDKFh+X6WCvS2kIdz0wtCPlNC58oen6DhIv3zpAnhLLfvCroDfQq1iwSHyXWCuUb7mCHPZ
rJbnFXTvBzESdAdwBj8zAPibYcs4p1uA8x2CUB25aqjnE/fVv09C4QnScs/jy68PLPD53fAo8a1Q
q2HGnFT0yTtdfpNjqi/UcJyiolh6ezQfREJYccW8MrxVKldWyTlU6pKynZZsRsDW8asxem53nCs/
PHUqn63+rxFeOUpel3hMV4+X1JP+5hohThEZ5fpBZ3V/SpTJEU+WxdkHU47+7U9npBPchWm5YAFL
zipmx0DoBCn0AFMWL/FMk0nijJ77Tmw1ZN/khvIeg2BImkkaNeuzBFAmim+uuhMJWPyvyYw6cQJO
MkVn2i4feiTNtrcwpXUA2vO0RHXX8POwzDJAfqbL51K83tgzKxID9s3ohiRq0Xx592OXDgC0ThtL
EXx3Haf0J/686b0i++ycjLduYyw7ZJ8zdTRVC3A6xBxPttuENPJ13jVVB++sLoFeg4OXYEDzVMuF
Tp9KWwOrJ40xjzPnvQckpEiAIm4jD8XLA/PgqOrdbzcMiVbRPaTvoS+1N/wb+JGJIgmZWgFbx1LN
vV7KlwuKI9cCSKoLXKnoYPbsi8dCmbiauqtuYCg8+/H6IoESLvTouJXMu+qcz7KQ6yiRlReBBCzx
NomqT3SJfdkcszLQ9CIl+/oCliNx58KfngXEQMR2bVxK2SLz4GkWNotszYtmuR5y339ofLTvOceH
HaKaBlmYgQSNIP4TMqCwiqtXHrSD04tHPsDsUvUmPFgpa1erkBtX7SEvAfMobZDCXv5va9gmiePr
6+R2o1mxHD8bSgcctU2Xz/gQ2qJ3pMpXyKNPjloKgRdyJuLDGW8Ovl95uy7Bn3URKfD0YhhwzSIp
SHRwqVdfiqsIh2DjQ9J83C/wXBCw2WPHhabndbYEMrtAAewOiRCSvKoM7mH8FvtDoBg8mUaLES59
W88lRG+pfylaOVq87OkMRFP7PvOiBHJ/DePCgHg+8LUehXvsq9Z/zMEc+ujseUWB7FWm2tLCr0nF
2PpXiYIJEjboU428AI3H1AJE17Cyd/EA4FNmL11wVHwRsDGey84GbV9Y5+VMoAwH7aJZnBbq1ng/
KJL0qR98JlyDGZ0riHBjY/k8eBT3PCqZSQElH9qlETgd95VVox7H8qbApbxmhaqdsswCmmhbUITH
v+6im2cyfM8UBEGbKdW+Y+w45EngZT0nH14hkFgHDIAUlg9RAUR0gGLjtIAhHomINO5nRnzztnvX
WQs3i+hz388vHygw/fHUSOfuBPM2+/Dk+HLWnv7Nh9LLF/xmSjc2BkDEfXjhA15m5yE6+cITwdvl
o1oDArBS6okFh6+nhFxA0IjP1kNuZDTt8l+Gpoa4ceDa4m+pFHK4o0z1OgrM2y5mZ0ar+eklmcP+
3Py6Zvv0ytpkzT3+d/ETOr3adOuTUAUHNC7ESP0j0zKzDNLZL0BxmOzMqfEbU3l97FMzOR9WAc6R
tXn/OzHohc24KhaLV6MdbDPUMCNP3y/wSnMpeZuC37Fc6VzI00kLzWnXB3UGNpg29BX1XaIov6kw
cNtEEr4pLugkTqWrsRlR8Oz7YggbxAgbXUu/+HT2oCpSdQHBXyxSATXUzKORHW1o6XR91ipFeZSo
ReZDhMVXz6U/PVSoMn9oSDNGGqta67f4p397EHbQTbWMnMYF99HIpEbBjC55M1Q8rZE0PhODgxPv
6FJYwo0lijFSPPucIJaD79RaDXyaW4jbdKkzulPXsptFON+sG3Sodzwe9M1//NNSTzgYfzlA1ROy
CXkiZ6Xqou9F/ar767glv1QTImGAfsqSgIZqdhhfzj7V9TxqA7qWVxOrBQq9kGJzGhdzCxOEpqj0
u6bhyAd5GsdVUxmKUC2GPR4YpCtsSVXpz72yVBglP7Zvh5jukGIzx80p2pejK3aNnuigFW5+ybkM
BkwC/CY2C0Wzl5r0lHRuUMOu+g/e/cc/d1nnli58C8opS5LXt3bT1QiIzuTs1oJPdOUJeOfyf8Bs
RwMH9hPe8+SWeypl2lIZ2X5tt2l5eC9/FOAO0maFLAfEOvbl8GyJKQJGNYfD6qSPRZjypP1gRh4r
o93MLp1lNKfRqg7gG1aoJ8n9+pSaQrL5kTKjqaJnRp5OtTmJTztzyrJr8+M74Ik0gYsQbuTCnqde
Wa8vQnFUYBHfnqounwfvPRMZ1S+yPgyPVlWuSZ1CdNmzf+NUe5SpmkeCAu/JH/uwR7499hqjPIwl
Dhn28tEu/N2ViY2ZrWquRt1LJwyb602aiudvDS24fdCVDpjfMZr7EOHec/7hPxZDIyzeVFBoftkC
14LuRaDepMY4tRtNAgveONEBIPqgqfALWaubXHzE8qBkNusdIxpZn+hNaSFW6Il32sizxeYT16Mu
QyDOGTQqWVbSCHIrCr0UYW/WAbAFasY4i0rSHuaOb5YaEdIUHSawTgDFyPNwhjFuuPbxJ8jieyPX
6djMRHupeKELlLpaC4WCVU8GzJGnXwUHpGbQ7I5m0TbXHRifetPW+6fO1TToRrtTJaINEWUc5PZz
NZbTp3phnkDfz66g4JxAbp4oDgfxaLSgFm2H7BhUfrHDgZDQZ0MnUXsV8JQBNxxRHWmDYt2fyk1C
S5fnrzsWXNceGdlikImsZ2dTjTkYo7/ANOtKM/JVfyNRnc8gGkqESBEVy3BnxsIuy/i5Qf7lkC5k
xj70/VrGEKu9vixi3I5eur85rtweDsU+D5th586mU7J71ynOGuAme+frIjv4qWIA+3PE/q0Y6+WH
ktvkwBdPqA4HfJ5Zxl7Sb6X0zwNuMuellTUzgeP29I84CYNYUFEwgX3iJuWcrz56C75QiO8hnJjX
ve9MCqbcw2HI3mWa6BKEU7y5sRjKD51HDC8zDRYTW+HNTJhHyNftS+AkuFn59tqkbHi1DygcP3cB
Z9mPe8LJqrmDxHhAHAbCeqKd9DQhfECqykczSGQoyeECQb0zNp0xXJH3O3EWT7CDFcTvK32HKpfA
jxcf9v7DEclH+coODGsALj74w9/sER+tPOtmFUsq5GNA2TlSQ/dp2UP6R8zVafJ1lq6PhM1TpQYY
2oaenXB4DlcqyYInzjlOTYQWawH94rceneAqpMaCw7zyqXSR1MSOyPityR87i/ooZTbpeie3M3tm
3wk61lNUQUqSaEsnJaA8hJMasEe+pB6UwNbIGm0HLl96yqrq/8UFXnHM2EE4hP3WTW7LcQVFjp4a
5JSVSJ1Ka7seXstH+bDTzKNsVp49WrPGM8EOok786wgFCk9E9CC2CFIe0QPetmxj0Jgh2JIRNQhE
vcawkzYupN0EucPK2ofJrZKBdFdSByyHJOxT+Q+3dp33sRX3B3BUginUnNe/F3dMENOVpJjWvchI
ap340PZZpHGCkfVPwD49/4pGzW2Lp3AQi2rX32BYtibgLNT+fhhur3y1nsxo1QiMQuxj9nDltfer
xf3K8uLhKUEJ5z/jAz07flCCse5fVe1eq28CmmXzIud6FPlglBHT3/t4mr3CmEKz0OPcJ1rH4x+y
Z5IILEi3XFKYOXitco/rfwCdHwEA/Z/a5WktXvGUMzbCNwTpPrafTY/lMmSElZlBfCjQY0bwVNsG
AAe4LVDGojrdgr9L8k2f4CteGBk3OkS0vI7hjjfPgWq69iRcJg4tgSA8MvH5LU2KXckOWnBvEZPb
PTANivvLH1J1NIJhg2LNa6RCsN5N7IxrXTKX3dakHmDl+ab9Tp/1GpadCsy5blCh447UDh75RWOM
wflOkupkNGYaWkpEd035+2LfYyrtm0jVS82Rpn2O73ib/E3twtq3GaJIn9kWouBu255/4YyAiE70
quFLQxGO4jU52quy/ZqN44qpehbSffeZOtLSGgYd1AclT5sOX7QI+lZNxFeGrXGkEVfmG+etIFJL
j+MRaMUGyvWCcNDvLtcNUcp6tSqLZa56O30TiLAXzdn3SOp7cLUg8CIzcKfW4qKe37nTdL1hQCNg
E0pi0E23Qn2OP7xR8lMrIPdkwj8ZUxRq3NwdXYcP3jWNXSxdSSoivSiIvqgQ2flkRYeykhbfInkn
AqXLlkptmqKdhYwXQ/lBZUlhWt9TiEtGAfLv91m+VZK5DcjKvZKk/bqCIwWhAfsvd2h+UL0ibqhz
PTCVxdJ69Rd1jz316nG4B7ReJQg04TXDAxcb4SBfR/6/sIJZKY6zRY5+INCJHLaIy4hOMVHSfutf
ylJe+1TWVqyWv2W7Gsw9xhCqBnuGmst9J3OTQABsBED9kvRLtb+xOzwv3OHGtrIwItPPIShtXxcx
aqoPCLFlCSE3S3hRrZhYsIMk4ijeDnA5uBNOhtlY58l+U00lOF4oeFLKcnJGvswJUAUa086tgbgd
X4jQWq1D23eVSVuLKMW8Z2yubp7Q90fsa9tlv7QX5zI7rZCXs5pmfeVO6jBAtNK5SVZyvIG1XTnL
3SVBv9P8MgcBPx02h29ZSnp4d6agdJsHRzFSSWiWzQiw4oeDp/+wj6lngcyUbuOjYtBmjJdV7SxD
MQ1voGElVJBBn6EQd5TNjQTkyH8JvTMQMYaelR+3trlzcF30bLpvApT3sXd0+HCOY00IAGjT05Zz
VXQpaJQaQfIGBkez0LSCJ+NYCluRZlnWUtBmJ/ktlxRfXnVawDGZO8FfkbpIXRI7dmZ2RltZc/fy
oFMZmx/L69Kj5tC25ERNqtRRWmye57oPJxp8NwiUk174XmGkp2TRMYFMU3kTs0dtpcl87w3tvLpb
96bbD3eqUglu6CggyE9+G+1paob/YPUDzNM2xLtwEM/6xtAr6iFUtVOSi+/cvuWZqByrko3PEAfZ
VxElJoFgRGCzTk8eP6QJiRQt6+RjixgrsV6Mxot0sfCyii5cprS+NxgRqEDnEsb4dXTFPDEp+/yI
nUH4KuFeJQEmNHe4Z9WvrQcXfdwWJev82nztgyv0/aEh12dYp6M1d7LNF43E6Qu9cqLa2/hnluEz
fVqIfbvrNbdkLR+FVM84iO4kEBhbaw3SrteWCQ2+g4sAiY7SbTghVGEO/yASdV9+lDzmZjfvtUdK
YhbEoxaZgZt1/mx4a9Q9dhBB5WanT6lbvY76Ehnlz+zE+Fdte7SGMvthqdSJyh+L1KY6ww76u29O
3h4R5DKTiBrDXzNYxw80n8cuePQ1U78bfd+s2c44YCuGduhxvz+tvO3KdjzaOZAYBUMZ009fRdvj
1WzJQohxgRJP63C2dlMZs5wUKFy5DTFOUg9lq/4F1IJSe5/SCmehQeyMZOezKEh+aIAkasN3e88k
wU+rNUQBBy2Rw6DK/gtYjSAd0o7++kpJ4GjII1o9+pMyLX20Iiy0LI5PAOWIJc4hyNRS4ZAkRFA9
o+IfazJpvMBJ7aApmv9KUf8Zim2L3052E/paz/9uHcgQB2Xw0U9HEAoiG0S7lPzxjtSD4outW4Di
7vTTi0G+eiLWL8Cw7CvswrXidlrGI6Q4XB/IseMjAFtw7yER5wHesPRt9oCpXSk1Ut/TGOEisSe3
q956lkkQ4/R2ISPJ2fzue8dE6hoWpSF40SSo6ZywCYNFHOP/ML0FYZHjFMMnLm5rRVEJuHL1xtmY
RVz3TyW9QoQrORcH8s0iyYmzH9VK5X2/anlvtxcbK5N/doEvLnYLp7QmMgMnfYd49jY7lKZidqc1
zIoazCjklayQehRLmY9xPPHD7zbeNohP84Ow7Bp1k98t9gJRj0QJm5wbOzFeqEkPgjOyVpuRKjOq
tIQKjSsoAEzm6Z20znc0dZsLsPfqJ4ZQQ7/SjZ44tRgJUS6dsmNfaXd2Oda2U3Pm9Agk/FV2/A/y
XjnMSOApH6KF0Fv1i+faZ5GtFYvv+MgMoOVZpoPOzjVOFGHpEL4GiFzogMc11gtoUnVfkwD4Av4S
8vGjNr/KTMTsFA/S3sjxKrmGz1cjgC0ajEzSr4RytaXhOOxZLF2vSMDsMNH6oTduBksRq2n4kSA1
xDRU3OD8VBhNdj25dlY8eI2lecTz/HLTCTXg1dzs/wmRWUCs/0fog9r4QTj3DIRlyJrv1z7+2XkT
TNpCApwckKdhBHXuvkrifnZhU0GsUo6OIpdHIOf6i9SnsuihPxP188YsuCacn0PWbzDyrfwbCFUV
qD91xx66QtzKGXwGX5CqZLLvRfZgZpNf0sk2oDm9sxaHEhnH5soASQXhVImi45S6VFdmfw9DYwEO
OJCTsGB5wawlPGL13k/qIPlLbi8gzM4JZqO66d4tcYxKSoHO52B86kuJTkQMf5mXw0Y6hs/qkkMK
QWigOxlS3Lc1LCVmgCed1K9l2ge6f4VtfzD2nZ9PwAYNLyoCHnZP8BruAgQAxjDuGzyYxxviF/D2
0OZroPssPEFmGP2j9KNSlJXzeaxA7kYgUiC5M1UoRr32NW3fpZGWL+ELqSdK1s1091PgTtKa7ye7
J+z6o5OfPfdAZWo48TmtecozIuZYRsMHM3lO2ykgqH0Hk6eQZeRH/yCqztrX0AxsyRXbrMgh5LPr
rFowq4VnyvafO75l+XzTrMBg9uOn2RPkJT46An2sSmyVQQPtvLd9x21TTuWHMS4MHm8XYaQty4JN
VKkFH732rGuXJadCbiP0IklA63DUoV32nRlBDmx093GqeZArdYx4pusuAirbYhC/njAbS0uoj/RI
l/+W+935Nr9JnMajdOqY3E0S+i5k65Bc13EwDhmz1VzyifmQZQTekduzn90HdKA+30fd5y/SloFQ
meBhaAs4kRAVluE1Nke3sqqbNS1A0SWwGyc0Z6ZFIAJA8RFRNi+ZycsDZkhfnLyh1eds5ouwQY5I
DqybCzejUJVRTwilrOtRmVs6/ccUB78dUHdEYPkIYJe8cQaIn3BjnMWUEKqLSfg9Gil7542nsAsY
TzOjdEmmREZtS0shj577YbcQ1TkiQVTvArAmywM0VRWH/5OJO0egWOFGvr8W3f8KKmhhz1KGcIpD
ZcXnWlHLix8OHrsT8mTR9Jcuo1+JFVS6bhDm6vfNTdSvMvSwu0jD96OU/vD/+yGcPh6fq5gPHSYz
2emiQPWkbtelpPKNX/eFrMrXWhS5xGaLaIkCoscVUBqexrR+MI5FOLckk4fdL3+3lgMRYA2o0zYo
5AYLaaK3got8CCaK9IxuM/rEftEHLZVXEDjjwX+aBTiVgZD3kbLtat6qKa+1mMKA5lDXq1tChh0h
w+xpc4BvPtCg8yVdt/JTN3tVQ4BxzxZWjfCSxS76R34RAc3wCjdbvb0+g0PI7znelno3chVzim1g
tx9IxN+YRJ5DhKuDYgslMc42iF5QXkrWax/GjkvaPJoQNSd6QaanTLK1/luIpdHEmeOXAPbVOgbs
U+2j23CbkGvdNcZc2czrwBAL+5blVRqLEUSl9D2N6C97MuM4Y7XZKKl1dOTCJVmfqDyAXq7eYpEt
cSZoM+aNuBZnz6W71mjkwjWtZm1g+ze3bZLgOQUbZOeArQ6iIiBgjfkawPQijq0BLJHw7UOgxX54
tZw/coI+O4muDiFRcHeR2JrJz6aCCvCeNHWxq2Q2xHllhsK5yFAJUj+Ddsy7QW+oqY30xIu9AEnm
4SGa16CIPDFBPwAm46qJoMiVtPDpmDEsBtNOL1VvLIZbZgwsQjC5uUEeOPk8ztl0/fwud/4ehmEJ
N9r2maRRRqJ6KeD5vcixy7H6IMjB2OBmmW0Adnii8boNiHV9QjjKbiOXAM+ETnQXxEEf2QMJ6Lzh
qLajZ6mC3mcwiG0/Dc7XUlLvUAZmvc69MKZ8MXr3UjsCxfK2OUM4J3Gm6HKnfTX+Eim3NAk9kmi9
5CCGzmr616/RGNgc9zDsmU4PI9Jww6WvuVZJNY9/DY6x+jaG8FZ+lo4U8hHnnwzscKZnTv8Uv8bC
iBlTKATfj1498FcEvG3vDpSMXEIXWYAYqznYO6dC8MJLNa2/NEUPphI5TrQPQr+rGO2RthcK8/0S
VFAAvEnUZ61FbTB2gLXRApyeRXNXLt00D6A2dyET122LHXEycmQ7dGICJPZXsAV2S2xzdZHXWvWd
Id0xb7+wNEkcwB7JENqVNBf3jZNbJ+cxbzNiF4030zQjKlFpNBX2Ei+th/WuuiqC4zZbg7xjNFm1
f4Sh8M2C0pK9pegn0rhdX/mOPmzcNw9ZQt2G8apnZLY5MZ4sbkUrhrwQcQeFjfUQMwmlgEtZg7Le
aUKudHohKFL8yxzOqQmyAzqjlfNizyQXKWooN5oNDbJYHI3lrhVDST+1a7SORroq9ne01CJkrb6o
c2BoCED/Xp4ir+DSqPomXrXgoej9IvJHmsKIgH/TQV4+hRuG1+MiagksHMCpMjvF2+Q6HZyHk0SQ
/brIFB1Ix+pPmaSJSkoYMoVjCNOxKd55AGPBTpEfXcic3uHSysQJiE1Yy1CCm9f1Hr4c7dJET6t+
mDLo6vOOZ+kaz3IvP+dJQ4sUVHRD6/vJ12MP5LJzzS5/xNss6uIYmwokAkmkQoO4hpIxj8keI/fK
YA+novz5DzywjU6A0CBhLtV6FNS5ZPdF42POimLdI2ICDdOXvYP6tIkYlKSyVfEAlHkB6N68EHFI
cS6fIgEE8gNo2AmD/OQkOiB2K7pmyNOCLmF+n+XhIJuk8O2R8P2Wflen2TmjxE6vIiHwWU4cyWU2
lb+Cs2zOPUPn2q9PUXJQ3JhfhBm8f++7xBhapn35UaFID9E7czKALJ/HjYOprjtuyDmMtCTwYs7k
IpCSxu6DUdCUm6+eTOHBQHZ6K8ojH5wqSESd+SdhNo5Mo6UoXyAN2kkEVh2TmZM/wP5OhEv+MnnG
WCo0jd642J2mVfw6e6hyJO3w1zyFpmJWzhpPm50UiF/Q5aCQ0B1Ba5Gyj6M4ZgZqc/VzvG6rU+t9
8B9eaG+W05nL7XZcMwKkscmXnYlSCU1XFj1CiuGjVicXwC3NjTylzPdKYLdqIak8Kg24EQWbu8sH
O1nLrvMRMVYdVV1hqjoXC1YHxw0+u21u+Wf7ai7XvUudsSCJroZ5ALidWxCplm8EXjVbityM96Z8
tLC/16+Pjvo2kLhaz2M29qjptx59sTLefkuXacBdxcmaTRODyRHmLYl5wZbOqVs5e9WEvQjjPii7
O6LX/sSgBF4E9ABTvg3c/iWM3qQrHO+d9H1zPQIASIM3KC4Yjutj9FKp1MIjI9kMkigrrAJaqD9q
LEEwEl7UiKaOdDkFn4DTP1UExchdMfzNTLFdx343zzfiv6DWsypTHEPw2Fi35tH4cI4Gitu6SzfB
9Ged61U/7s7KAwrcSJqtfeVTOcr+mkzTIVcfPcBEuwIb9YTDEl+zQpIo5MtY+PxCEwOAfmBN3M9t
H8NGW0TjLWYBQ1wAS/Gq6ZXJPqwq8VNfmMPvOktjGUc1YAZed9hRduDV/X3ZXOXGwI9iXXBJUk2m
4uPrJn0XK/I2E8A5ALHHKisN47GPYvpMWhUw698Og4XQRtSmbluNSyCZ+h+x5Hbrt4GYstGYRe4K
tiJpXoJymUl1yQrLXc0pZ2n5zXckWlMv179tJOHITijCgSA7Fd/wAKRV7y2NDEParxqVgPGY5JhL
VXNgfA7VjA7yjR7DIWh8wG96WMROz8PePxu3+ChJ7x/qLVc7ROaCYwMwaVNDmC60F6pXVbMi0EXq
ocydnd6qEM5mkva/la+J9I6HfV5k9QoHsGErNadfj3ukHbG92/ZZtjvaL1RifO/Od3RvCXx+SN7V
ti1SQh0kjflon5rflsZsDjVaM50WvfCjfQszy/B794QbYH3ABNMI/TTejG5L4UlCwInSQ+Hs2R+K
faylKij8vjRbaL/Qb/ZPXraHgfCN6nSmanukpC9BnHSU99Lpwol7U+xvGN8CySC4GRALTL00c3ed
u0v+juzJyVJJC9YGIup01dO7mFtgx6Kd9J9jsmTS7SJoDDHvZeB3ShbNtjPfwSxlP8HvEWGzLEE2
tH0m2Cn/2++HFPOnKbAB+oV8+IneuFUfNPRaRSOQrfWSaMjF9mKYXHOhJCxwrSd7woBth7CaT0qd
I7aicuZXf8EeBqoQSBDb6jH+QkhwfuJhQBVlKYterEOesEfqbtCKXE5VFHRwWkVb9QzQG/sAfOEg
YUDAOuZDpJIZ4OSQBZZEFa/NZPOBLmpim9gEbb9KpqwElhFVMTp/J32X9m0pyPG0CvSt+75rC22Y
3t8ZriIhKXx8VtbhfMg83VWBmRBy2lx7n/9FQTabtDr4zovP2LBANil1xg7xjbWpetUt2YmKWOl7
ZCjykXToo0Vg3woRxK03lrDw4glNcroiVSaKrfzFOFolIfwXfg8iyHYvNyFFHCjsQVktfvsXR88c
a/UnjVBNO7i8zmOQv7f+O/R5LRPEcnCMKu9B6lF/SdySVw3ComeNrpznaHWgxOPf9ptn/nZXhV+4
seke4sz19kiDSUr4nBhWJ43QRdaeGytKuc26gJ4lHBYHzZWhk2dUGrBdvLqyEJa68Ogd1NvA47a4
vgeaWGbDfy9W/eRPTRbCR+pf6GBotK+FAQZsdpwlSwWAiN244YEpeOvc1o4NYuFtvIQyQIi+/xtA
OVC6bfuz7JLH8C6+eQdUSgusJ/JehcjLxe1RajDPRUbCTh9N+4RdbhYfpe4Tz8H89hg7kgRCMAb1
XAC2FCtWST9iyRl9zBDLVoGe/NjbmSOC85dDVidVomt9ze/d05rYCwrunf4mZTOdthPCDBDbwSxE
diwb6p5/jyS28XnfDt9yyvxkr0yH8N0rfCOEs5z5gMGF3nWHSyFNucndgTW3HcCauygKDirraZkT
PgNBsYyP4CAZ1u/QtuFp+eG4vFZftZF7saFKwbJxwaNoCcNeWAznbu4Jg1Bi1zxAvcX7ULBZ4nwA
GpD2sUzGKF8UCv+NtKTXCdmi74AvAP9IrVZFQyLZtKrudgOnuBki6XfRPMMzsyFfAqJDIoMiVUmU
agIC0kpjPGkgv7/IqZlO359iulhmhvMIJVENMwFGSPeXpJ0nd8Gy64kZNLbT54MScXKO2lKUDryw
QAa3Xkf5hiOXy1t6Oxd4X+KvBHeZEyA/7kFPHLTboHtcZqzt599FLSYIfv3O2U8NuHOAVGt5XXxb
MEI3BkCHjPp0h2x3/qgCZWZXqlAU6sxMSCFfak535SW7Jp0OkdIz+nqSr0IJzI11JHvpY1x4/hFS
l6iPOBW6AW94bcmJnl0JdlsW5wbGzTVWbLez+8LTcbauaJt/ULbR/e6wm/iqEaFVhJA5qjpK8LfW
dhAKC2Jvf+135Fb3RbdsEYwZgQGlxSlflpbbxhm4Qi3F86GBm6kpfvuCSQGAh60LwhNtgBXUV8Wu
/S/U53aeXK6rm6A/cjd+0gtyrcuDZBcqIxap0V7TzatTN40Dm1UXmD+k+o3dY9xZkv9JpIGxh6Py
gXV6tWizzcAp/5x3uFGp9oJznsJe++xj6iOtpK02V2wW7RkjXsaF1OzkBSSRu9wuGrbClV0MUSft
wwc8IbKPLcDMq5q0i/jpN59fEu3w/jtKh85HClI7t/Am7/As9Z1HKc4e1DRiZtanMpoWnxNxBMUj
XXsUs4zOUwppTB9ZxemFTLqLXAnGrHJdE7HWd5X21VbTPcFUBhRqW3FJyZZnFVhaGRLVtr2bFbR5
L+akLbl8AA0+0p3WY32BvQzEeg6tE9WsPiK6a6BFYVxswaFaqFNVulQA74H2/InTf4qbFGrg5x2W
elWp23Ak12h9mzre0/GCWy8PM46z815z4HxsvyeLMB6qfePQdyRX+LD0QfxyfDR5KfOVrUXgt4PQ
TTK4fq4O/S2TMsSYg9fHkItuctTb5WG0Bc86zY/qZrjF1+Y4A8gpTdJ2P1hMK7tiJHxuFUQTyFK2
ZhGeqNHR/sWoH6bXuvkehmnljtJpUkFxfz9C64JexZ1z3eFxSRYpF7nKirTXIxn8+TKdtSbjowXs
PcTLlCcgXII0PbCR/be75ApFMPhK1aqWAAwPdx8GObTLoV7bJDJEjNjJ+nzJxlDh6ECC3yhgfnrZ
aryZGUl1QNH43IYcIoTPiFPfE7J6W9LtZoXkMqm3c9EjePdoBjPQOhjliirhnsi8mboJZkgmWLrY
lyZ+TpJVL770zHzW/D6QAgTHdN5YdaTdfqOWQ9K88ya+Z9P623S2OLQSkTp266jd+8h7qX2VP2Bl
n3CSvqGTNnRlu1q3za17dmjmqtUaDxYIJ4j7bIosVqseWcNmGwzCGgcSt1G5rHKY/Y0HFpxAqvsF
x+2W/ceTgnAlip7wAaHfoyMu7GuYLYe5b+LO3AtoQO5XFcqzKFCdKxkGTE/9ODGp7Y4CYK3bmYFC
DX2GyLP5JKAzwUojPmGEozObnMN/9nzaiSJa9ESTlyu6YOw1sWyRqHnCx9wLCbuTwMXUj7BtbyeT
9IL7Wo2RspD2GjI6BLJFaTpC5az5XNsINsCYn6vWQZb/5AieseUEKRQpyb5WJnd5JGdHQ+4iQSxN
Pg8wEJRfuwhsIRZHY4Iyx9not+Cyp8jRdAUagyUF/oX62QV33D6ck7qy1pPj4vJpkcPV452kXToU
3gXKdJGdmpepyoiMce1pOGM5j3iaocb9J3tocfik3H3pt6QXiaSlnr1eVKIqOy+AJciFvIoNs37X
V2Z40txuCFYn1SLQXyU0UIaV82W6T6+Z1vRsJdqrsd+i5voDgD/djkzM5VQ+n8+qaDBriorT6hPq
Lj/SocFPpgJN/k9A1x7IRIGfW+Yq009hXypFX+cKxwiZD7+VnJ8fkHxBw4w7LNNfqdP7M/1YI34D
WtVWFAp6k7gfy/h43lLCgOo38PEtmYRZa409P0C1+FpkKvSBywaRa2sdgQ5/GW1t4qXz+GckicKN
3HzOoCdPf81SBL3oq3t17Lv3Y9WMAuse84XRZF9nE0umhvUTJBhpo5utiCryT6rry/ou8OJhmbPv
HisKRabnbZMvAGEzZPA5BC5X9lDslSSVR13PYAVNba3Wnzt4z6DYjE2z5nSabxs30B2QqjlszFP/
wzBZ/7YqMfLbUXCdZBtzAiy+5GMBtGYWJRZgkCIxMJOKv5j0+/PlvS2pQ75iqYjkl8q7rlBjI7js
KTfmbej1XO1Kf4MKIOv9yezUCt1qZMuvhH6l4PjLdPkVE+hzmriWHU89MllisfPTHWGDiPGxW9rh
UwMB7CtCLNyW6d8BhYmttn/arMYGvtRo9PKLxPPgPplTOtniiWKXyyp/zs2d7Oxf1JsPCXCiUwo0
AM8rtAFwmqIp3rmQVVfPytqyA9HhvA355o/RqjFe57scdc6ELkvR7mmLPMIHG62I+tVwZijITe2N
UfTm+lfgNBzBRSxGApKf2tWRK3hpDf47628oVOUjyB29FMbhQy3e8Q3RSCLJwSYHN37UOkSqAytv
iNT2fMwNAthxA5m86m8Ne4gIssauFrx39VnPVMXWsiZLQFd1k171jbrmnPJuVlTPt69IlZA5noFY
HpZHDFFXrVQTPK0irHk7oS60pMmufK806xx/YX7XAaYdaYQuUuKr2JvVA8hgHbazrcRuW6+Rb/hS
ys0cIhLn+gpPvGc9YwTU4ZQ5m4pN6Zwzqx+7HCgCdCnkq8Gi3wW15fkq9FWF/FG6Z+bG8yL1RB+k
y9k/qEsV31EspbPpThkzUlNcBLq91v8S6yw8X+vfR2cGTkD12OMOWMEbCE9AUy4OmK7yejA8V9cg
l/C7+NtcM6fZOJBQucss8/sq+6MOxxh3ZvJsLo0HA0OZnOnUVQq10Pl3xmlA9eDQfzQho7iQgkQW
W53JyNwGKq7pa1x/kA2wohIdE/hCNsI8c5BIWeTzsMza6cpQ5K2+rhd/nQq39Kz4xq6QYX7NiyPj
7b5V/Prdw6HQmrxKRmi31+DYYiH4rUgGkWHEG7EFpplVfw85Ga1g/Sk7yOiDzvZNIK89WDKjeo5c
nKVUD8LQQ7MTSYXOxQcNXelAMOXxfxVFldA6wP8qpGyprN85rtEFxqfRFyiUWRKQ/4skR5phu9nw
Rc67s82vAdSxRorzyicmqbEQcPU0PkfOII6Ea718yArhwrMNhSiaTe7GfqISOs73e3j/URfKYD3m
HUr+LywsncDk5ljxYUc/6YQqaca8LTF05sN6rRQKWJtAvIfGRfiwFqqtePnXkgUFmVp2BHZmJL/S
5sihG5u/5Fu0aBPmXPw4nbckKN6TBKru7lIOqNxQuPa+rSUUtefhsUXvCTxF9LrHdJIWyZ0PBcRP
RSa9wo/n8tdhXLYUzXRwF53acqJR7hx9myO47RV9UUwcdmMNSv3Yb3HbjGiDscSentEWqufKnYX/
8y988ptKqLLdLclJGPv6KtB+rRaOW/29KcXIRbcWF/v3k0cFMYiK4FNx9gbbYxQoicEY0Xs1WYyt
+O8wle2Fn63fGY/6i4Z+hEuhUoybPi/naJkBYSue4ZcxZ1suu7ef6ZgLOCaw8OZsAjexKSkVIyra
41Yk10YkksOK5h/wl0bjXhj0mmnMBLLVKWcVmWhwBk80YGgPAA+3dr1XMHDCpbHfPkzbrLC/K/uw
nVjO4GpxN3idLsUWYtxj0v8dZzta3MJPaKx9+50kRQBx8TTg6dAwu/2shO4qBeZN8GR+eWu6PqxU
3VWZQpvS7DTZMIv14i45PAphfWilEITyPTEB1QFWiP2ENWQqA6CHmwjxiEyXh0mwdXbdy4moBVo1
JdmguOM9S9kuFd7z+pXhX8uEKYr/eOhfgyJQtLI/GgnCO9VAqjaz5mxx9niJD1DIEQ8+cMch16xp
ehnTfj7hH37ayRm1Iw2b0N07WlscDZExMh3JYSXnTwVOdeYL0UgCVbKovCGjmU/Go+VWvb8yuzRy
iQjsA4E4ZtP1ZVyCBJ/e4P3Ax+mCVsr3EHwwpJGmBDhzs3J32LfFvuKQTXoWZoG4zFTbrvAHAlmr
PQfmWGeDDfIIXFoyWCfhULu6SvPvQyXgKcdhuEozpHx2ynAGq8159D2INhx9PgpRYPa4DUTDcsfB
R5Bopjgt/yPJzdPSjwD6Ndte/u3/oVXB4nyKsyAEkbZHxK6TLGN6DRiH84ZeU34uqK30lyi0idhm
bBb+L+vRk6WrR26vCbcw6oWJWnol5zrgJc3yoZtSd9wu6uNo3TWvWri4SC4t/C96zd7H6QWytVHg
/lz8tS6C527rR3/32Ak1FuBmtTrrkfrZMAyWWHUWlGEi9Zj4NnRC7Xkezkr0KtBpcFZL5srmeYwG
ma8pCezqoGVmoHlwZeys9M4edfoEcbnCiT/iREnuOI+asUYKbhBCePEQFYGNvbRH+zsZGUBB7Tn5
DfMVoCrymX2WRIGywcD53WaL5CzDj9osvxwVgb3xCHJYgsLmBAJwi7ykkeUdg1xhVEAZUbc2MGfS
OJJpsKgiI7A3FB0btZm0ZqpvYdBWgeq8+t13DFHCRLmHZ0Bg4TOJPqxF1yqFHTyWQAlKwl8gydAI
w82tprGY6nGzIBxiBECfIdXimXKX2JNu9gy/FvfZyirU/DWAxsM/IoO1C7V/QxYZva8OFttnBjYC
2MF8panDfzdnvWI36hFv8j0Jq+RVcl8cjh23rKR1zIo3NU9o3vU9snXjAcgacXjrCy5GEtlHiV3N
pvaTtmRZq6O87xcKsd5r3HdaXuWfT0vcxnazobIP48P/cBMMT8oNTDQ+vObtGJWGL6fl2muAKDKF
mQ2F8VAssQ3c2Ffbosj7gdddXSi87a32v6XMmH1aRINNsWqWxTewskxW6uOoXsPeUR6+gr8dix8r
WpuBBLKAE9pV7ZiKvVJIb8l0QsZTl+JP52S+8gfvNDzZ5A8EbHV1ID2ZC66J3vXTLnFwXpDnPK0A
j+fGGAdlPahJxivR5aK4+ObcJ4Xr3962gUzIl9XxxAY6HRjBEDQxwATwd2omPreXRpqS+JieDutA
aCoyYpk3Pdyq4UbkBI+0VGLNREJr2IbqN89b/lbWrpCMRpLElXhJnqSjaO8hF1VAgdp3sj+HARC7
lJUra1rF63hdvYV8b9AvjWzTK/v/fmN2s/433knDr6+2L8+eM05fBZeC18q7oRRpiDrFKw3f9wNT
AI7ZQ7MT2DK8ikBLuJCReS+vW69/q+eNaw8oIOeKNQnazBNybTqLbB31M7ZoT0vrgsFKcNP/DgZy
OLJDRAIo0hqPVuxdTX23XHoCWZ8eKQ8C+JtHHD9pSLz82L7ZdpOUQ5XdkClb4o4nS9dLnWCE9+L5
nwr+B86CWwXSppio5bulOEdz2DqOankf8HZsnjriMPtJ1k8sjQzwGsGj6j3vATxn2foc4BzWT2ZG
9fqmnN9+GWSN0NHnlm+OXt/omOAjfdFxGwLysZeX2aA7MG/9TGkggGCVUizu4WMQS716GtsbL+Uk
722I81NYUtCZBn3Cu8BxAx18QBmcIjErY1Awh6mslhad1RMQfMlfO2xM2js2Q1QmkE1Wg/fbnroY
VrCiBNvneTJgCN3NJ9TViBd5kBMmte091UQrr83v+Aw5yNOTqWY3TVQe2jdEpp8NVlEpWedrlrEs
cr9H2UMQGnqWequw23iQsuqvNHx/6s3TeTU/SU9KyL1P/vTtOfj6ZCSx/7d77EnIzb+74NCkYYd5
ak3ICZoi7pMdob9uOZ3wjAoXFA3DpFQGgFFNcnKq2vg0d5+Cd+yGAxEwrpDUiLceFEqG5cirQNq0
vBjmuasZlY1p1ttW3D3pyhMj9wSkRoXsD5eR5KUMoeFrQt4E9KH0s3P0EgiCxXnEnRE8PmLLmmkV
JgQivcM7vJS+7cAThe/IqBXh4/ogBTg/2tYkJQ56em6rq5ivSf2s7ZvheCOlPprY8J8GwQxmwP3F
QBx5jAzAwrx2yCAqsvdGLt2evaZJ3rhq/fAjanJ/u9GqfAKvqSYnI1CeFFU+4UY3TCmn2QOcfxRZ
BB31tvUVVKMfnB0FT09ucbvGbYtms5h1R+EHZ6P00yF9GZjIFuhKF1mFpX1ADfoUuaj5mw+5I8aL
nub4NauI0PL16wyjd3y62JAszHpa2fu+eccqeG5fk0pcsFZs/PAfU2Zq7PDJXyCJII9kK2SDvzp/
yueeD5zOQpdI10N3s6oZ4fwqZ/tfvisfEr65TRJvU6z9SBqVhy9ONhaI5Qgx25BsDHRGFRpSwF0S
Ky+SDGkOQZf/ECdBpkeGsr5Bu1tsO7/1tCx2uh0YEygBIb6xQroUB/DnH79LZHC1g0ua/yCII0uV
KxCh6c/xZUsnDW/A6F4DmAEthoPFI25F7/CmeNmI1YT+mY70GDOYvPQO8rqNHHVoiYiMwqPvf4Qd
JLimgVV7DrQH74AvuCW9DYicKBfj1eE2UIg/h4+rqmekKllzgiVO33o+Th9Z8UfmfpYty5f8lW/0
UrjaarONQf1vgKd3NYvp6nuGmj/UNfvSHOUZJ2YHcZglgRRFDlVbHC1KPG/DGwB9VKTUusgTxjHo
ovwMYkgdIJboRjxqU4HJQfNW+pKRcQ6ByFVI/2Wiv1Ip+woadEZQUSyZ3hngv089f7AULu3ea3H/
HrwgYnDhCTCydOOUXo4+S/q/ic2ZuqzGzY94uCNk7kNd3x/7G8hipEGV59zAFpCYWDQLFFDgWtXF
YiGsPkJEjV5SyCrGjhuGp/szx+H32grQQkrj4LO2l9XqJDdfDmekOLtPpPo54EMe/Ojz8uqo2o1c
pZyAk6CObDfc69thtpKN2XJpwnOCP8edG/qdlbPDlaTYwYBZZHQiabDimo6/YSjJ4iU2yaS7dKTX
gnecoB7+El0fHBPsbiCQ/9ijxnCjoA7YIcnv4uA4RF/p6XXEHWiO2qn9vlk8vfPkQAyIVju9DXMz
xcYP8Nx2akfbog29vHiExr2fjkUzphZ/Vk+HhbFTicLEROQNpMm5bn6sHdHAWy8I7YY7EHCMhMT/
EjLr/W51Yz0cBKcCHZTv4aVpD4aDiBVDCI7G3GeqdPjysaVWwNjQ97D4g8yNYOcLg8zhxM4HwgR0
6M0uB7S31qUMfTk5wmbC4AtQfOE14rvfV+TvLxQS1l2MEPYHOPoR920X0HAmMKjl0FwWF+BzEW9Q
hbbeIH4RuMPidCgPXi8OgcVGJBQ96UPA5Pon3HWkg5mIMfdfhn084VP5vst2i8J/myfc724Bbtnm
7opIYFLjr+Ld4wz/Y/Zyc1yCzQAniH5/q2kxCjKTCLlgHNb79X9W9rjOGI8TRf2I/PTFetkgBrXV
V8XdI4Vojmze8qgcHtQpLvSMkw1gBoyKelJ6iNk8Ppbto/61PoEe4jUx25Jcux/pgaiAZHSFbJpX
8hw8SISY2EAUXmPKcxkP+FU2lzI8O0i3cE5LXxS4hGX+zyEGFbPVrjukO54MFiXoTfmnV8M4A9S2
KBDWm5StuZfC+a5RYDKWreMRFkL86tWUTshsHKG2WFqjLiPuauuZ/BW1tuE16i2XZgrrAD/KQcFF
rcsrK8NagvmTbnhofg/o+ffcRioks1M9qFBHzBureYXvzyPrZntg4WFYOBilj5THiGt2s2DyYpZ1
KJgs52TUv8ngSUipGrx5G39+MbwQhcF2zY5pvVDUXlzWIBMmL3sjTV1DllpQLwMT3wzau1xt3TEz
h+WkFlGnk6GlA9fe8Ddn5U9m9PJrlmTRVNAwJ2zXHRcPAlMtzRa83LD2hT/mYRh4PE7CnHSRokL5
BwcAlVj4fVzRvadbS0gXqxLEgz4ciqLFWbhju2S2MOd3ttrnYBBmhikGutObI22djvV9GuTRT8hl
iZZY++dMKOtuhq4cxQmke7947JIzeB1KbN+Yx8GWKO8jaIii76gDpP+EFYHDysPYz3cHWrfx2g7S
8fPp9CJvgJJOeY3B42HwU0GXVPZrY34M0QEWGqs2L5RQ3+iyoeg5LkVdwH5iALw1r8qYGIUDQgfV
Y1VXkxCrRwZYttj5vcUeI5VdaCl6n3+oEK8yLECuNcSnUPgyh1g/uq2panSzzWbjBEJdV3MOQ8ge
6JVEKbbhsPYLVRtOfcX18ggfMr35P9vdJR4Rj+xZVNxJNb0Yx1W5s7q/CtxTi0GZf5tRWmyKeCXb
ey4smbauxkrschs+4qiITGikPT+/nPQBQ0DD7sioFVEWrNjU1iekmAcN5imR/424zSKOS8h9Vywv
rKmPbQFnwWNQvRDDsD8lL+Y97m06f8oQyEwUxa/bioqHnxlfPaVuKB+7+thEb6xXWy2JEonovTSa
mvgPT0eKJ2xOAOXUntvsw2pGaxYEmpQXavWYSMOGp14q9lOM0SXGf3optCn8SmgkDhpn6liJzBXl
KpuSC0YYT35OxxL1oKF2yVuCH/lxInA9tIZviTcn0+xULPLKiWGVMRQg3wzF/CNh17Q8xO/7U2EE
7fARD4iUzH4IMOldspFdZX0msmFJax0qx/wLutOhwt2/2ulK0Rg8qGAk1b1rZmMBS+Zep0XvxnmZ
slqWI99MbeNOYcGgINKLLaFTvP8wVaX2hlVfQPrVse5B8HUNf4qMW0W+ECTCImhSM4ICSkq4CNIf
5o07hsEKCkIdz97cKVagN8ZQCMStlKjDd042N6KNqkAvgc1UNUqdy9GuKLKFV/KW6jh8DpohWP6g
Ypu2tc7VESufz+g/lJ6kiWxgxU5apo21a/UQI31+rbtiJM5BtUS4t8DxfenyhYLo/K/3w6YPUo+u
A1GQlncHDxfwwZH8eRQ/wdet45ql1rU4xZb7momyH6T+VGnTNefmgT2kEiiPB1fwAkqcfQGb4oyH
uLkKtWMTawMGMehH3TgfdgVAkM7JsV8rurV8HQUpeAGuB1mqXmQh3Sz7JVGnDbTNosxyZluMZwV+
GQfsZcE4l1cVrVwe6KKvAnNWzImzeJ1QL2glkKqmhzv3lSQecu4Clm2g2YwHcD21XjSroiy+xwBf
kp2+koDUJa8ZZaKdG4TIfVpkURPSeONOKZpsTFnyTIcmWOFEv3aGcb/WhjW+AqgA2fWTEArF1coi
wo2lTOTJmgCN2TDM+8IQ5kk5MQbcH8AI9Eip1fxCrF1wgQicptpZVPlHEJ5ZA/fvnetkXOE+NEiF
RJrC1eW865GAeK9JSOuTBYJC7LNDbnrg75AlMVJPdjgHW6EmvneqVLfilJCq7ztV8fed+jryTit7
taQveDswbA+zBQHk3uTQn1nes4vHbqHyTbHqcqiTbPnWwPtMMhYMkIABJOqaSeog7cx+S11CIrxD
FkWMBJCV2Sr71kTZqs/dI77nmxhx2hJrFhG7ZFQQakdkK4j5FMYOWaBBYBXggwONx2y9l9NgMwV2
oubrqfAsbj0CL0h9lyOMB39zCp5odtm26P6fQshAb47ejAY7kATPhXwXcwJFyIOq0O/gOMpy9CjB
8NhiaCJ2vlq7qKXWilcCG5FTNlJ2rMtptwTOqDLAGNS8GtUIYwjPAQVRyChpUm9ZbRya5Hl0r4Z5
GOfvefSttME4nMJ10vXeHefNU4EDITo1PH72sxnBBeybcwVRtjyIZ6gWKvxt1i17LDmzbBHnlRMc
SP2UXWd6kJTq87kbF2SFPNlPpshIcxpdFlanWxv+x/N3416/2imHeLSUs6XZY5nX+JtvYXv8zS7Q
8pdK3nO0vee/SW2NF7PAWNuzYoI0U39bO6pqV4bqXnzooOpp2JVuF8mYcnC3rIJBrl0U3ZGYyhfI
YvGADC/w2pJUvoTdmB4pMF9UVpeOh5L2ExW5fNkCUTUFUKpGKigEKPDBHN75bj2vTRLn5dogFDd1
AwHH+35ITdGHbGpY3d7brbAFvB1iXpGVnxcxxdRU0kfT9itYkSetqr19Nqe2hzfGdLF11g9TKHnl
FSMc0jjVlGJBd9zxBDSxxgzz8OBWhqi3c0q2KA5tdU6pRYbPABWCJAUmogiK0MLiciEBBkakQZ6w
Oyu5z1WLQlrMQhDmLlPp90jqMQmwtGV1WnPrWfSU3krg+X+Xm+wKy0TLd1JuMzRL9r7bWXD+2jCZ
cxjHj/8sQtKUoRS0AChLLpJX7K6pNEAPMELJ2rjC1JNQLzef0gwtdk1qFXuBrLFA6K563xkO1K77
PaVpe4ltK9VU5gZDe5pG4n9fmJj7CkeMM/dE8+cJf7XLoqS60+JLXjV8BL7FziFObl965Gtd39EL
DUYmZ/k1ivvXrn//zouXycq+s+gKnjguwrodiYFOVOswhxhBbIsR4WR/PhOV8TYTArv1IR8FLIRg
Eps3HLcjTblYo4BGJQRBJue1R2YsL7ka2eHz80I6jWL1y4KBmhHfTSVJsOMwHKr4IWxkdpxB239E
IttEJ4enFd/r3RyS4D1440XkqmhfTJ55w3R2uvaL6zQjMWiOKjgGBxD66lkrVcYAeEnfpsgqT7t2
10W8CKEnUn3wM4ddFAnQSI5Q1VkyLrsA3Rkg3G5h7buASoFATRtTP0Sc1VodDLWwJwgJ+Xl/eIHN
ordjlHJjZeX0qjTyvaOwDl4jlXL64V6FwWrK+lvKNQ/j35n1zAXIgSyr+RFK7wy0rtM00imAV5u9
+9qWPMCx3KtP8Y8JeuiFVbzV18UagNRjbATcIfgRXIoOfbC05ffZOmql3iCbN9yEaIOK9/oMlDWm
7fl7IQ/ZeJM1DjxanrSOmjY8/jJ6eFztPvqcLtHdHr8SaR6Bj45oNll025oG0INpxQ5FcI315X0X
szzBfOhJ8A5Rd/1MuDj2OEuUprJA4uTzOBds+ZFsdm8byc1ESyr1aaBunka8oGvToueSchoAM1Q2
QCd6ZZ/2i5wga1LQBvX1PIJxQUDnjuHRenXo2v25mKpfaFAe5sEaPsLVXrB3AS0Opn08WvES4G6y
fFVyNXvKdTayskRG6mdNAMYdHMNYY5yGYz6waZPh674YJvlnIerf21KhgfPdZdmg8mux+oXP7cmZ
T2Ao+effeF/fiAFJdOh6dXXLA2JZVo3zXZLbRMZ9a7xy/VJPqWQeIbHP+BSdhTxrfWuX5u7yCsvj
DlJqHMXhGUT9tiUrBcUTXplwF3qljDw+vIPXsbkbmxRfKQec8r/NGgBdeQBByySFVmPPuQsfehvi
df41WVHwZp+Dyyp0BkNwoaeqP8L4/c/SxKDJSnutGe7zFEfaX3eKHMoZdnuAKYHNd6TtL61UuvB/
cbzngsdHN/XNG6OT9ZvN9iUnf05WmTcn+EzQh5wv8X72+ntNXVVbTNXbtsyuP/QwiRPzQ0YRBrXi
6nzZ0pVuelzAzgkf3vFjcYCBQu40qo5V9/gjPSCnFjFSX5ug6joLHXMv5YAKbe+RQB16FTtAAQZc
ryLveI0dLiAg3FramGIZ7Lzj7dYAuwJ3nrVdeJM62icLK/pnkRSoAd+I66YFs/1O/ntlWMgcjAJQ
9qs+B68JL56mvDtglSJpKFfrmxrfUWp2LTi5z1A1UMXnVu5hsGS6UfTI+4sG7gRtYsjpULV8+Nep
tAnA4xGZjBbQK9X9W/yTNyCjLKCUcC6at80FOxsHWS1V06Roaxg7Z8J9txvyHZt45UB3fwDmysrU
7oz0ZGATSnUlaSyEPekwz17hFTr3bgwT7yfyKvPX3FLKbYU56RJlAaz3eON0kjecc7oh/iC41Z/a
bZ+UsbJNijzBhFMojNY6kqd0180fSKzjWU+O7ZPVHOlmrjlNlBVmH8lZFoaVQCNpYHoPp/YwLtKx
fZjJOzDZvQ5hHH2vP6EMZq1nK/xl/n5XYI3VNFdoSkLfUXHhjph3jyqd0cC0+cIHq2YVizjUC+vL
bCJfXfH1m5xESCej6GM0z1SNlYE0MC2Bl5of0lOHbwiFbhPQzPBD44930wg3UEOd1goiXmKWIYl4
nKhJLiorEpsLGPH2syeUb4dpUHREHEXHXyqGpUrOmxWvToo+n+XFtCUYYp7ETX8dCnXoA6JqxHtY
radIoZ3GOw6rRyqS89hcxKbrriH/0JlCgDp3PshmWPg03xRAgGeI/XZjvu3bEBwPhZzzacGwHv4V
7UCQkDP0yOfVehQ13UuZPE/Srd3k71Q0qnqew8Llrva62bXwxkNd2Piy600zUCGV07pGVQQs8ef/
WWbYiwQ+Zhl/qL20R2NpeNeZPvyw1F7OD0rBpOEKwpsQJI3CRSuF5X74ICAg9EAJh8RN7KtElmV8
t8q7PC15sCeYrs0YYpSm7pIrjosznCA6t5WBJAZRg5XezuKPRuAGzIfOxQbEUxtm0QjeXJO0Ilf+
OkeotX5LxmtDdAULxg5LUovgvYwT7soCLy4ENd/PrT9Z4DEYQLqOgSWe8alL/msOBvqkl7WR548x
HlqR5s84XvTT8P47fPbbvyYmrXylISoq7C1UvvT3aQ2EXQyYCoVLB7bBBNCrQU2aseXC78nER8vE
AhL3ciiwv/zMrPcukfc4pcBaZmBIgfTRIca5MRFWYwJ/LSnzuEcUcB66t/R4scfOhMZgPE68AZSa
tYZH/UCvK5Ojx6pFZ6ntPHsnYGKLjhj2R7iIF5nacQtlXrvK3R5VM9TjwABPCKJRLtDKGVVN3oPb
dEKFb+jAh0bfOn2D8vQ99LSI0b8X1Z+5HrY2cuz1MQ55WYg+I7OlFRBrvasJM+oayVPr76obed2O
dOk5jwkm8PTn7rHg41syELHrArjrXc8dIJMUTBM4p6q/XYlJND8Sb2gJ7zKxPI0MSvqwHD2X+S4g
lOl2Tvm5T1qWQCoROgBjb4ENujVRnAZy1navBV4AZzjrOmCjg9QYcohkQpfiLwJDzqzqWpF1Mu/e
/hdWlTcn50fdR5x4YgH2PSdf+apM3nYRqSXqlTNmoXEZkOT8YI/ciz0+1qybLejNxM5CvqX6q3/8
41IwlatL9YQJfDKd8TorGb/1rm1KixVYDdiIQaFDFMwvW2DCIY5CWyzw9czCsYuI8hzfwp/XWE7h
W3ZY3MyMo6Vm17A4NPCRpNhCfvSJj06DVpcPELTnEdgmFE+7omGSImz5l91+8xcXPKHZjO3KRt4S
1tw0k8j0wZygT/RB4MUG/kRL/iTn0WVNqqFRn74yHCR0pP1TYsEhIlqPHr4ebJ/RQlbkMh7dJT72
b4vI9ocOf+HA9Rvb4QIjUj/p92qVpQMf2kRabXILl5PV9kdjR7AC/JQkUqkud3EUy7h1RXoLSrv1
nK9Dg6QEoXh0iuI1TErQqSBSFmQCkvjgjV6JLQtuFoBK4YzMgqCNYt5NrT3h4GDLn/SgGajvddVY
/FJK7P7K12xUOXeMSyegTs+qnyv3Vnwn26a4C6dTP80r8PcwALcRu9oUJHP1VO61fBQadlpfvr0K
7aDEV+h5gczQEnBWsOmMnbSth4lj68y2jYFihxy/97jPTbuzSNcHgGrgCxoP9heNO0/4LVqy5Qri
K1CkhLO3VO4JH7h4Jf317oBGyxHe7E3UPRzcGs/DIozeeS1kAOClFlesDhyKn21suOecl6RJ8CZ6
Eiu4rhzm9WyOn6+i+egGQr5PZZ62/7Bc2DyEQQEikbrXo1ppZJYh5YRRjtn/qKC6IYfXMh/2dmX2
guzgi5q5gVg8bmpxHCbNGKLp/BZi9k+sH9427d7gnadLaqgSG7Gijj0xDS+2I8tcJYaEBvyxFdZs
uW4eqibGmJknp63iXx8dA/MqOiADM6iHBKBqsJdgZb/ESvwA04Utw+MKZzvZ1knSiQpoLFS7K97X
RokJwCzQUSs+RRZ17MlIFmSmA0LRgFoM1b611Pw4svjpoJkhhkY+V2AGHOQRfyX8DeOxWnBGET0q
KUstEyL7Y2iDA7Dh7bH/YGsPNqOqtRhJ1M6BNyo7cGMXAFExHS7ETOhAByvyVrQV0ql4AZf3bcvc
xXwDQugsdae6AfJE9FAgIJYPNZRGE/WQVvhL7+3uZGBg1yRAdR9TIM7W+KNFIOvhFjWSiqOjKdEZ
g5cnrkyW3N6nENlTODn3KlQLJG647hJnLzeukjlCAT4bpIWIIxVRb7grtgVJT7QE2aZzzLXo/P2p
ifJDq+PkSWw4M3CYp1GbYw68pkw409lg1Hvh8C/sOO+TyFbd5F3ggndjP22jdYRX1hMxSZT9f1ju
JbKXbwcd01oIDWr/K+mTZ5ua7nGoZCAvHMrXPIPzaUt/TcQqrQpiw36DTBq/qA9mAUODV6Y/CyGY
0rAzPORXEN08gBSQHOqhF95XUx2mLhpM9UEQkyqyslBS4HAfXR8DJ/JsbgBt512OR88uADg4DhvX
l/A7Mb8TwDA7Eg9bEhjuctuL3O/qwRaIHUws/F5f7hp3WrTY8g+p5zOsOvqSVxnmjKRlsUWuVPH4
B+8YkTBw9XbTEUyXoIX9VV0pAxBx0wQGi7UkeVIuJc5Fzz9EiVhpW07N7/OKF3+sNp4eU8zC6E8G
783/YIn/yFoWqWKo3g27xowsXT0G4lsRr51Kxpzc0Wl88ynRmLBjTXogSIwB04ez6nsNNC6sW1PK
GwPvDXCEEG5WF4WRqoNqnxjdBHqOFXDzFyQfOIsK76iDlBVqmLBl850OJwkmth7UiRbJUdjBQl06
jUbF40AneTHd7PUPbiF2Yc7ZRNR8kf63yjfqcEpVYP2rosJWNGXeN6y7QGyamTvn+ZL2ut/uTjoW
XqG4n6/bjHWI8VnxOQmizbWqtA62FdRtJT0/MTjjAJXPvcM9L4zpkjfVJwXn3ZhOV8Hq21shXQ9O
jdSsAWAswa+20sRblC+IiMovHlrS4W8+CAjjnN0rDalLfsvpJEbULPeZhXsmvQFHRlIpV9bQmia0
MdetQ5YXDHV1MkHJilpAH0aitCCRsmUKivCeh0IKF3uG729RhQDQzwgyYN8E6oZZ7IAePNbT8xDg
R1eG+i3sdA5/QEvfgb5PeE5dzxqwjrSavTPXuBweEjeKrCNJ0Tvnj/D3/lVQZliZsOU9RzRuLA21
A65TBkt8UmxVXcooUOM2QVOLVRVD7K13ULgu2FFSAGxgGdke4Ryp9CdTaPemb/HyzVGAiIPSvnX1
Be1auhoirUWqXslfTw4p1pz5/H/kG/6KXUltut1OtFmFj7SLNwhm82xa1KnzZMGjkyfsBPIzKvrK
QAyC+FvH4CCbHapoMvF3/bOq3MuVICyLJLW44nbtIbMMg9c2E3yfKtQT7zlcHssnJcot+RMjjTVj
RYsID/B1niDJt+yotqQNDslldHIJfU2KIXOeWc250v931I0aUskkndjmw8wGd5YJOLFuNWpT5boa
Lcthk+nXZAKtZHb4uuJBAtt4xoJMeDCBGRlAXMtbU6BrV/56zdUp/hTbUaw7fnFpvc4EWf9Ugj9y
P8/MlmGNMizWxfTrLCFG5oSO1i/MiBDC8sM0IYDeXq1F19MLu0in3tCmN1QkDwV7xyeZhXmD1XAw
7dXl1Y0f9h/qHgiuAU/YWY5OYCsso5uyyQG5bDnYCzOi2/dKTDjeONzgSWXKw4JOWXXuO3UQ7N2a
1KKf18hl9Z8MVQxY3oW2q+03sKUFN8zZeFz2C2XG46WMOYuKcT9D4MfXn1yW7SlI+xkBm4OSYz2C
UF+JVMGDz2nlxhBrZNJ2DI6NU/Gi+NIEws1xYYNj7NLCh8xFNqr/VlumUDKisUqUhdU68j7MnhEy
BU6X+BpVOmLXyx9+ZgrZlFlA1osykANuFu+EYibanHhVsOgzVMQw7hC6v26NXdhkklQwcKrm/xdU
EohOv7v9MUTt+4hdpdQUh3FT6L48JudETTdMdzvJzsdQnEy3mMj54CjzncDk+Zt3MJXKw0YjbBTX
UQnGdK915wGR613HUOW01e3EIqDkTx7gVD29CrbHWyjcJxI6KJ3d0fmmBfsJwQN5aUtjWScSM9Dj
r6M1DgyvsjcfUA6/soCBqwOaL7kt6onN68VzRBzi4CyCaydlB7a9xdeVenE/Ya2Ud2kHgIWIFEjT
zxrwa8qiFSdrXhrhwF4MvXdaTKOnvtifpj14hiwNtqSLuJ8tnEs/A3f+2KjsxJPNpEktKzepjej9
+w8PQqjWOkxQEUcZvVPT5ekKVkK7r0K5CKk2hszB71ONyeZ0BlMk7MVSNf7A+BdSGdeHavvfgCeB
wIL0czDpPCBI4c+E2k2CijcYYsu4m1ys0XeKsNchk9LXNMOxCgBtxzn50f6bqQ+xt0YDIZPKIt/5
0hwfn1yyLJA2OHlCva28bpaI2vXipGfiw25qMdP06+iLsek3UrglhEDV5GlyooQkPMh+Q3+ejaTB
xmlQToPOCQe/BJDN21ewQN7PQ1QnNUpv0prsMq9LCavYmAfYgghyRHzU8xVEcq4sl/GaglpIeNAA
kMR9Yvbs8UOBKItpn+f3UxGJZLeBufMsyDaewJljzndTRLNbHl8+Ev9nsUgLUHlDSMWLHY8v6+Br
W5b6nwg5GKSt9BEaYXmOEr9fp+vO0qjsP9i7Huqy7/emdUC6hqIrD38QPBwL29hjSpWyGxv3bBI+
F/xatBjOcVl+eaOOGWDLoUCGf9DUT2nHBoHdxp6dCEydmosv5MqBL7tR97EGb1mTsfLIJn+ouDK9
Wj17tMNMsLffv3KSJEFabWLcQwhLPSlFgc5wILPuEXDg0hy+SC+Kk1+eu9qmkeWvUv+0GvKcZhA9
Vs6ZzmwAWpFKu7R28JZCekTJQF/2QWJJFeyUF1KO+w3SqFS0NSSvwtwUhdAyWbND7JUo9i147O+G
aEGG0RIPRQvPDA+vtb3C5bO4u6sUDbkKtKjWont5+7hgEci3ZveeTuNJs2yKYBX2QJeh/aV6NdvM
eJlaoJEVyOGYQfiuUGXig6odylVWSqs5/wxAolUNgmTn0BlJx24I0eQ7b0i+lJ/WpU7S4vg4ZSI/
qb5kJ4NiBOQyMej/CGO7SZMjZugjqaPZJ7nI1eI8lzI/f8oMtFMCwTLvXy2JKp9Znm3mz0Y2+S2Y
2qcMR48dKK9GOU792wuD3Y5LOqtan9sVrbtfV8xcJn+qEatWPT19u2jx8dNL1pngrW8VwvFoU3Z/
Fmj+hRpFCPWAxbXg6NBpmCP9seRcjkXIlaiKBOiMooP3OSo82x7OwGtunvPbiFO1rBseccKYEk8G
D7opkAqsEZJ2tIe/yvGQBZy5BqKPIdQvxY8RAsu6zh4BPd32Za2dFprLyaAKFVi8HMZDczbXcjBU
JZYZ0Q+mWGkDap1dqFX3wCxiEJO2I3+ZE0mQYAOpv8a/hVr94+KbBD7XFZ3OQ6/m2hY6RuTLE0AW
KVXu5fdy9lrb6SmeGafExH+S7FxYFkWQwzsn2PLj0HhRgUmIOX6OEi/X2m3uD9v3OH7oOaUy/mFA
pNcOj3DKtR+uyOtLvm/f2nX8XLR51Z6B+OuDt96zTpqzIZtgdemGrTU/CWz1UNrxKOLoW1pS+Omq
KCGq39+BIoCzNFFG1GDt/3ytsUE6/BfQxDGq7vbIXfrIY4s9EPaK/Ya+XJuBWJ3C2niNo9ny2b+I
AUMQJ13uJMnsbFeoTPmnyewSAAp5SWOvjZg9SZNuoNhsLJJN9ZUaJwhHFrTY/KzGYiZk+bvmWjNW
ov8m9NI1nFXK/ENIP/c+Gla1GOvlcmJOiZZf81JGZpb/H4bbAykeeVfgsrpVm4cjHHM2V4NVWyLh
/+54tmDLUIIFJ07wpVobU+3lypaw8notg5tS48N21iRHO9i4fZdHKchQAkf+VOsuBHCxfmVS2akQ
jO2AEXhpzvjuNgxtUAI6dLLCbE3fTpp3r2+/06sfRAlxN/vDqJXobEA23NODwkXHrOuSdV786Sfo
hXjGG8xTFMiN5+lkm0Jb0+FCny7KGlSK01pINkQKvxXOs1vTJ8GIG8H5yB0pAdmGfPTWlnyV/rKS
+oB4TSt244SLYXer8Bi5HcHz9Cr4NrYMSp1r9yURPD/f3HcnWP9MGr5K5Pb/j7CcimZZE+OC5ach
BQgv1KEfBasIiFWd+2otf6c8uA0yu8alTsAKYHsizAQhp78rAMaqNo3/ftoQC/7nlEHL7bBpghPp
YqMawJXAXLpjpo8NWIGhYKlGMKy204+/JM92UpXlqe9vWJHlAlDeYEcqo4GqrXjJOIGkOKtAh1Xh
wpHkS8DGsjCAdj3t36ZQZMp6pfCZJ8UwJ/bScdNzfEFXWXId3wN+Igwoo73TZ3hQdNubpnGGJrVU
6OzqRgmvXHMA1BRzVRCp3uM4OxNTdUrV5mRhb3QRjGF4nm3+DxI+MiM08uluZsZ9JML6tMk0++kr
VnZjfnKsQwOYWy4WLDRtjrss5BxorHj50ePsKPV1Hrrmf0jNKRtDxkkIMEC0WIH3G6SHidodjuOC
p76+38NDoUdq+2aiM+cFOyOmblsyBadlMqgJVSdIzBp6fx4I6gnmXOcZxIyQEgCG73dNHDirIYKE
DpJRNymGsSWeqoIcFDkRO6kNKMkk75zVNqXpDUuL0fx4YrhKNB+iwUzTx4hhDrYrha0ooz7CO1zZ
nS4Zbo3G6sMcdCHkcQ5OgxhiNbopxnY4GOk1lQ3HmAYZoJket6PET4cBBqC1+GlChXPCItTpE+nm
8GRyjfmB/hCQ7mkMv/sRIZa7T57MJnarm0mPHFk/MnKip9e1TQA+Tuv1pSWquPvs8lCxUG0QSGAA
ywelEVKfnboZPDolmtGUO2Qn8CBNMkUoBAe4bN7kmC5MvQeP/6pMUs83EamP/iHw9u5DtPLiWyZS
w4Q56EJ8RADc89ngIyTtJVnPzoah0ynBN1AysXe1NZJc9xf+ePjPd1JWbEdK8qdCAbYtpy3KTCWz
RaZSCxwBzNlC1v8VSCoyngOy+tOqL//97xXn43E/LbgjF8LFVBskDTa7BUTbZo/3h0+RZ0qJBAg5
NT/XPjtSo2z4aqi1+K24E6Q6ju2OCOrCw2h8x09RhouG0rFC0pByDvD+VXzVOgcx0vQJQUpqeCMa
iS8jrb5N9dNBHY4sY/8YoMP+oyRziPFjHgykufBbnnLuXnsPrXpZYrG8aGFYNZL6y69/W9BnFsP7
CjHy0Wa/os0LGmvCrYhg6jXkgelGIdYwgqU7xBjgniusZ2/7yXRK9EzyfiPvRGlPevtl/nBxNdEz
65jVcOlVMH5lWcPVe0sIFkEAPSCW0twtv45vDyXti+66eGlFeAzqmv7CwS/sIuM6lCXa5yr0Q4Lx
ly5EO9a6u4Ne0vlqAOQ8+h4ROsjj13qL4slkAzDk3kVY7sFlzFLAxj0lS5Zr00G7p9iAhRtf7bHY
DN40eqaruTWtYTDYiljz/1Rj1tsq+x44M40K2Yal2AVwuZxCS4CF3fRDuy1jLjNvW00l/zYx/LUV
/skKtA0chNJ5Ui3WrZVQyOyGnvmNRr8YGsnfldfIEu7nEj1641pAPJ8dFoRIppG3N7O3yMX5fYk4
c/Cqd4Vg0JrKqYRbnsjfmGtRY4e18kaiW9EhNr8S16cgI+YTxKnuTMWl7HuvjrflFJ5PFi0cBNQ+
NEMco+ilem/L57/k+Q5OucN45JWu5+psGOMh9G/UzImsS1NhQaxFHW+QhiZMsz97rx/nrHgsAQDs
a1njvrBM8bUX0eBHOkKzEzhysEHi28h4kAP0H6FCmmOl9ogZfqVbXmh6fGQGfcQCmwvdI1DSZgUd
qVQiVKn6wiVjZgPiFeyBwh0AsJJ5AfFdK6TG0ExFbOmJZFs47vJT2gEHgwy37qBQ/XYA+WoKEnr6
Zw2hPlpcXc8hf7667sr+LYovf98aeSbt1v4/wuW8fzF74HyfT+aaE2Ug5xchLLwnxfFZ4TNse+2X
WvDfH2Vbx08JwBrq07te6ufFQfoKEKs19m6AQ2335EPkYQ37HQGZ5tT/XajZY5GZBTMHlvIzo9z/
2FsDrFdUSNWHdWv9Ffk15iqVCjuQJRd6vLJCpfBpFldXe1YzilKFMXD3LQ6E2DIprLa6AgCOa1MY
uZ+RNKFlPiMLL5wcz7dX2GPyt3dEyKKOdhC8S1EMF+fp3XRMuOSbPQ/oxn8FGJ5+HVmzvSZ8CdUE
37+5nWsEFGLnop1wv38TreM20wyowWt4sZ91Cj5a27j2JalPkpE0OgjpXx9CrLZr1ExWtGt63v3U
iohgvnbfMKyaMsRwZXRSjeR9GqImecY99+80HLSKSV3TOSdnfvWUmyHVv4vVUtdlsZvWYJcA55dO
IktXNtK5pxjm+Nbz0Mr0Jii4/o02FSlpcDX8rF+TpVIlQcVRBvw0Ykl62UbFp9vQJ0P0x+NFnJa4
Ut6Y5dfv1+TyjVtyVWu7OEtfgeLS3WZ2fn6qdokHpPs5UFdjp5JrL38eO7nIbxIJhlClPfBMIP+H
hEZru9goEH06Kg67IcL0Ng1FFf64S4i/AAnH95vnWmXOCCcuQ52+wv91uum+Hpj9+UYQrB3JQxli
cLRlyKo13Pso3qlU6TMILKjgA/lFuu47Lknq6sXUW07YmOM93/0f54tLwsX/maJbLMyN6DwJDhe1
WtI1NbwQE9FLdFbzI30tdlU80DIHfgFAUkWkes9x1v6OBr2XRuchyR81eznh3G2ilZQWXCoteF1Z
XV3yvh8/rd0nDPx88ccqsjGxDEX4trAx22UcqNeCwDpetfCDl8w39kXgv8pDWWWbfMCe/jQ+aW/h
YfZKhol4owqHRO/d5u+uqXK9KFMjN7SZFZVc34bYl9ip6yCDwkw2dBkJwbvkImirJ+gPe2JgNPgo
zjSZpzYBFePPNfcksAdeC7nMCt4gEDntlw4Yq5dpkWQB3b/zJpIweIs2bQ7t07ojePGdAyn1pFxx
94Rus3qsIY41QJDcnPFNWrndYoboPsW016T9GR0/eorj277NjbcmR5pqQQQVh65pLgC/mNdqTW4x
gyB8R0myta85UopPaDi2yZZ1nIYHXsjuEJ/99k5alD0PBXP+QfbbWPuLE6RlWauNFzxTraxlczWr
VKQZiLLHO1mQfmlfXrVd2+RAsy2TfG0FGqv9qYTQyPu4ueis8vSPOtZtMoT2u8SPda1x9Tn+dVD+
MCEtgBWkbl66Ca8/FMfWT8dYSyK5TgBL6ejY7EBbE39HUf+Pld3woXbgsyoUvwuohfjH9o4RzD7p
ULELixX3ivYc+QiOffMQdJDcIxxESd2K7bjbSbXdzE0Cd+54i5ezPTJf1fRyheQOn6+t3AevW7gO
xscazgx6uLcw2x9mvybHTcx4L3dZRTX4QhZGVfza3R8rUy2dT7GnbiDx1jL98wCz4Z/yF4kmmxKJ
jrFvhpkRKLDzEnplApCYJs+SiAffK0YVHY1w6tGi+7gzyQPi6uAMCV32WKY5Ykt3L55xms6UUHTC
YpOUG6Iw7SQTtQKlfqN7qQG4+UizYA/ZbnH4NfX4LcBbuBmxBRCWauT08p/6XE3THAySjRIb1K1j
AGlNJAot35TFPEsK2Xn5f4Ju5ng+6P1ms0cnk0LCKgwba5pp8i3L4gSNHTkrhVCAPnzM94aPCY8g
3o2UVyI7zsFm1dAfhc6oK2oDIZTcm/8A/hp/vjzfIJ03cYRlCXinKsMjlkvS2Y9fNusBHM9696Gh
P94TmytZahbkDWSj9i3TwEWw4EISpyQ3MlOOaFU+P8ZxAL5gv+vU2r1L2/5nDdprkjrGlSt1Hp2r
sSozPR3q9eZ6luVqLNQ6KE08U7ArYk1EJBCuvoHQQTs5ozOapYtDLiZL8OBF9KybRYpP3rtBS6m2
V7N4lv2Mg1oY5FRVbt6PfaYTNwOh4dYP8ojdLjUg3hT488lAc4GaAuN5p9WtwL/oi60C2USHx/Jb
SdtmfQ/e6rm8iKgdMbQRNFuK41twcnNGAolosxQKaBXvFiik3ULs3Mut7I8PvYy/CMeaKeOtQ1vw
98kV7G20EBQdRGBpvAc2Tqp3MSZinprp2r6h+QrdV3OSqlGF4RrIG1eOCQTAN44dH7J8gMt6SmGS
410yqSsBmGohzgthq5/WoymUn898LVRT4P3pNCfo5DAV7uhkHk4JBOgLKAytMQayzfTMFMfQITrv
uCJrWZk0kYMp8ijDU+z+0L0Patwa0iFj8/ByMMHBbiCIIY6ITUPXHnvXbQHuevC4PGdNuMwFxpIj
Abubno8JOhjGwA7+Wn3KkSkMTD6HFDu3I3lN51N5yQPBvfnm+Qhc1Z0K0I320jigZj7AAhYih6zi
OOvW0Y79P2+8z2HKFgmAceqJdk8OzmXaLqdwJkePa/HlS6qEHf3r47Kj1UGGW1DolgCNOsBE8LNK
JHeNXAqAEUDSlPZjSpy4nLJLpYwZ0IDPQwrEidRRp7KoH1YgOsXoCXfHUDhoEzbwVLJNIhbS2/2C
WtsMtl5wTcOzSn7oxb9YuKADfKO+/XHo63BkxMet9IibyrvyzhZf5JW/7IVF3g2WvClg3AXdEmwl
9F/C8VguDzu1NEwN+xs5nBDBgxHUO/nJhMjzVjfiv1UNyFhjuBgfFhtFId+lFttamoAi+Ta8HfWl
N2oy5hzS6m5AMCa/H8IyRpelYzTznecsq8x1SoJRQm5LtnR+ANoyYapBObd2kSjG+kxMuwnpMqP4
EewyXVa1bETgWggc9qAIHwa8zjjL6uT6PcQ1tFuC2P1Z2+xtfg84fizFNfL2tGfanF3Yz1lRmSlR
aq2SiOlc4wN5EzgIzyvwVL/SchD02GLPtKQ10LtwBegMrful8u4LKMwZx6NZ4rVjIY17rqTLUzUW
RFYIGq5VUId3lT1uahV5aFEsdVD3/AHcFXuFjpLe/nAnNlxG61CR6FD+Y2Z+tTnLaT5F/zEbbcVn
trRDYxRhqQBVciOzg2MP37GyDWGfWEycL5m6wp2a0hO9lmKPjPXUuSxZJLpVGPWT4DDK/uhtHkKh
K1t2GTfgokayOEhLYWfSlpuqZ/Vl4cxJn2IanZIkRJ305Wn2pbGBKxCl7IFyTFJZTFw0OlIOCU4r
po2DUoEGJrf0CwPl4PpFaWvLmpNYU0y6dRcEyWwRp6BSRoSrFNalv8yeligSsxxEyGoAMiz7D4uR
HzzDv5mf7VWoH+HnhA0/spoDbnwFEM5zSC90lU+dYhTJvwtGd428OnLg2TQdmeyUemdXd1GdkAgN
eXdQvNpntXoHfNwfpwesqv09eCPB2hxNhRpDco9qxaofHYO0m1qZv28xjFK3S3YD09ywrodRE9Nj
0alBL/+quIFDEh6XPw8r34xPj8ldDZiFlHrEwbActJsBbUOGShl47AepxlZsaLZAX1VvkSXmXdEp
OZmPSVvlIm4CuI5gAkm5nYG8+2Aa97Bq4ef+WZJY7hpUSNzK/3MAnC0abqQKhd2t3f6QdIbuPIiT
ywafcL14axQhO28+BppFl6mbiZ0bTQfIDtb8zxi4AFU+E3Qqjh9E4RkbN4ltvdxpV/pGbHGsfu1k
DajmQEQhknaEABm+IGVgay4IA47rGx5zmsJ4PGYQ4ji2FS0CdaTRA2MvWe44+bAiOCCsCDzwzhBL
hY2Ms9SB+PQwYMzk0huF2MGvKTj6MKaYwc3VWzZtEwBW2S9ntZTAvnLewFNB7QWDnMtRhdc6q2RK
fDa0qBQH9YbkNidpVlnY6lJklQ0ADGKhuk1bxGDEs2LnYmu2omVwyXP3vUBp9rfDRg80LhFyyG4S
81Q8stS3tAppvxkdhiVz695hMTmkkMYqAP0plaolCY0Z/1r7FeUW8bhgFheWwVtqKv/y0ZwWUS+4
fXuW26UrusVPHQlSxrSpDrEr5Z3yoOXLkO6DJUnKSUZHuKCNx9G2DsU0+tTg88mcYATYrMXaDjJ1
Nkgs0aei8kn06jEPbexfvmpXPxEAcxOZIVnjvLcHMYXJ6tfmsNqxxgbrCNt2Oz5q86wm8q43B0JC
36hLLtnJ/SCN3Owe0hGF2pj1BjAh5MyRhkA0AKg5cNEcf7z4W51rZBjZ23VJ7hXeWZ4tKkyRhXHz
jthNoaOhIxPCza3390PrWQ0X0pKI63KGDgLpxMKwKwpdaJAwIvsm9Z14C04591jawOJuYRFlmwF4
ViP1X7q0iaENPJnWuUd61lN6Hc7SKAn1RDsZylz2XbqoOTKrrnZe8AtNPTRGzzwSesyyb0lHvj7j
fsnXCB3LFlquyhjwgUZj8jQ8g2pJgGrC3EObE4H/Oxi8l4Ii5X+TubEvSRYUCMkpclrjjM1oYmlv
9NQyLrkYruSfNTyVcc8uPygZBMwzk9U4EOkMARidTBwMMSheTBM6YhYjp/6HACK0s4QeRyAKBGOA
Jx2yItVMFs4dNsrgQQ373Mx9mEqJ+XegnNR9K+M9w0/9i7gOzqCPYjP8d4Zi5fRKStyaOg9C4xIQ
nEfgoR+Nm4s5GLpQd/8ubJk4+HJXrHngdL39TRM3h4Uq1VfOASUwUNpeckH+gLL4Lt51pxk5D5CQ
MY4EZ6Xgoyf8i+74isGAK/xvIqutGwGl6lSn/sqMv1Dq1IjO8k6nzYkXht56FyJOm/Bk6I5FwuV5
88K2ngBCQnt7yyqFEluxVZR3gVB9sYskIc90kLZUTEArPW0VCNDrI38DlPTDMHoj4uEOlvGCsloN
OmA0RbvOHDnZp9UVcHubb1od2rKnHcWqpH/MtSCExj/HpYPzyAFZluZMb18+2UQcjtd+sQ3ZoIoA
sSkJmbn4m1osHcDpflbn1g0FlTdf8fpCw0WICfRXfkmvYBA6VDaHkJjaOhoyr1CqTt0m1vhth6iQ
CoD5C9/0BR+ZoAqurVM09xiSu2h5vFXN73tESBLuRZ7uuAemMJ1nSl1TLV3NTmml26NcMZfE7jpt
EJAahDqGHO3ji6PJr7t7ELXHaCH8kzKNwXiSOZLJhxwWKMETMVFmROJSrO2R/PDJKiEjmTE80hjO
0OsGrmLKmTV6S/668WcOZb68PWPf69USGnCF2zlg6triU3JntlbZmxuwggK1i1uefcHlnYyIH6/F
6Eo7AaNQBegzGHNFIX65JrYTskOxJyymQpijnLN8W6fkG0ZvHVtnD85krI0zoUslbilzZphpu4nN
cJoAyJl3vYWNktvWF2D/3gZkjg4TBU44Zo27CyOeKqSKzVAW8pnWc3JLVITf/yZRJBZYvYRu9yc1
OJpvcTsZJxqgs1woAlvO/GSXQ/+T2Ao/FKqeArKIZ8bPVqjFkNgM43YjPnr0jN3mYBhSMtETwVT/
f/eOqSbX+e40okBHE40K+EsDf1gFpM8trNj4Fhwvzpe7t8aKyL3AxvihXYAs0X+CESGA9ggCRv6L
eHdhhnbIAXVRot+TOG01lRq4nOFDDjCptNw8tEZtS3Xf/k9aQd9kc2RGOGdqNmpUlyVNEvT4nKUL
ZBWpGX3AefmjRF57sjHvku+Pvvlo+z3YLgHz0Wwp0WdEQgOtzgglxGW+ArxhZSYzD6EsZxao+FGA
DdNwLJHV0owh/W+32yrtMjulDLUFcL6LmEtm5TyEmXmZP5ecNlDyvfBgeXVVdsZwRwDEkJ+sg+zg
tj8r//7y+g48qTod2jWnYbSIqtaW/ba7vCvnVU5jj0vwH/JSWIgS27d6P1KC8SAKGyB7hS+EVker
0Ammrrb4C/Dwd3bNXxvuWNbhdvZq2iMl7ehDBAA4Z3tPMnzkCTaiG5H3zX46HCWRtYXF1YrFtJEY
6TNA2JzCM7clobPJpk4Av4fWZVJ0yA+q4hHoCQgD1+qKlbdlLSjIOHGQ2virABtSbmqwRlk0CJua
S5PLD/NKA2vUK/tIlj8nqqB3O2I4ZNibiSfbcq3DRYp/RwEnQ/zuOXe5n/62fXhUxS+OSfOafkoB
6eQoS7cX4BiocIg0PWiTgnQALsIxwQCnczU54lqYXr7b+ULV9ZnvfDrTT66WzFvyGJXFuWJxaSV2
WDeyVz7CNF7c1Zei/2ViEB3Fa7rG3H0WSlQJLUjJuH9TmKHFXA5VQJv9XWNvVnyApRE4rIGUzrfj
Tyz8eYANx9KD2KC2JT7rtWGwgEaW4XLS3Sq+Qo6+qyNwR7JglTpuYAYt9hHZRief9LDVTPCtyBPH
vk4s0RSyGm7PTGtQC8BNbsVF8A6fWxJADmQA0AJg4lcyeRaYGgRF+abiIwiVbaxMqT5NTxYW9cCI
b0u/c44/0dV3R7hRO9aMybG27dOzgstzZ8iNKtN06dem9SxSIFXMCjCB5HbAFKweOKsLT4VY8TvU
L3Y08VN94eanr0CRXr3mZFk2LJ7HZeDg1x4EKfHu55Di96ZaeP6x6bKYBJkc1JXL3lplPPDFV3U7
A9mvgQE/p4BJe2CTQ3q7+aGCn1VyNopX3wedNkYbDYlWczrvwJ2YoddSIXK66VetJARV8CvLNeV9
HYaeLfFAfompHZELXmXl/sqsp6ZGKqrK9qPXttslkNNe4SNClUto/UnNwEV8Ov6H7suYC3iyDV7n
T16nZy8dsAjI8m06P20b1/Js7ntXKkn7BXAvz+MYRIS/pKxJa8F8MoDt5idqZ5cq3DeE7w1A0udy
HOYd1tNEGZLwp0VzNZ2oBV18rxulbZi8WT8HLJvI+SWlA6Bqqr/o5uOBGAA8Fh2N3g+ofw18WZxT
TEFeDQhyBigZH2dRaabTnS3IuMNEZQsNNEQ733osBzwJVYnAJ+61Ypm9IMwKhtJY1MOpCY+z48jz
sJ8JU7GBs8hMTIjtistsFzIa3ZQF5DDtN1rt34X0r7TbOqn8BY41JbjJmMtLpzH0JSjlZNvKo2a7
jeYeFGIxLaaC3RyxFDe/4cPC7o3c7QzTEBYT6PgFmoiVDy+ipTy5Sl8tGV+J8jqcplU+CivIeItW
FKSL4eXuqCEcQhZcc3RIrfxMtQR4g6u6xFeuhH5BTB1U2zHlj4Ed2Xg9MrYNcABh5iL3xlsQFuXG
0wHLjvRpGH2FLlnP+UejWvrn6YtCSp56V7x6kp8zoz7IX8CY9oQCFoAXaAxao9QDwq+ZKFtcBO9F
/HYwL9qX5KuMFw8Cnm2o4unMBxWFJ06gOOMFoLnWIEpQVtCFplcV1Tsose5rkiU+rSHNCZ2l06kN
71dpb4eYKLjwgiXR3pyduoc6F1EPTmBllRCVg5PJj2MtlNwyEz0KY7inCNcg54Tq4lxoJldlGf2Y
3ksYKHE5IYjcGxWJFFm1xVKQdMBMRQED47ucVR+EUqKAeLzGwDG55bIMVRH9kDBLgtz7zF/4a9Zs
a1e8Ae01DEkj1BQXoIiXQm298vpf0D/Vu/WInzuXQL9QPin4pU7+OZ85FGQUyEHI/GBOdjGwzIMB
8iVioE/B7BwVUXDoliz9W/KBRpH5QsbhTt+0WDbu/kAilw6PdqIDKHJFrFsOxCez412h8PTpz55K
1KinxoCQeLhDl/PDtznJ4kBG30vN+mQH0cpUVxvW+3zaWXMqhQ4RBoJouJaSdwqkYbeY0C/T7ZXM
xxKqX8oZ6XGYhUMIE8yRV4N+PfIuJV04lLFbQtlNcj6rP5sBCbNlenTNAcOT3Yf/ncDnoL0NBEjZ
VKCHg+iztP4a7sS81P3yPPxMGo+3hEk3f3B4Aqxs6jzwnki9SUz6f6C86SXUm3AssWcHcwMpX+St
JABXlwhhGMjL8ySyp3Fiy17t+sk5GDYiPnB44lCxqLyAn6hsgpeyu/fmo2UNpGDVIt8gGVmRFKl3
ji3mmueqw6b5u0PvvcPg0eZWabyl+fqg5IJ7oi1t/+I5E47hElZnXwn8XtXThleMRpJ67e/Lrqzh
Nk9LyFDqWYCb/ZDRzzR3k3EyV/SgEmkrmz/xzB1RAJWM2XA/M8GzdX3gNcA74fPN6PXlA5HqY9Jc
KrRnifGr4Uz+szR3vDScMweFx9QAO8cLagfe6iatv7Bf6cfaQfrtePl6qCzPnQrG5FHNO75pLr5R
6xlpdFf4k3Fz8UExCRP5r1IS8IAMOVz5yBrVC5vJxQlMmUKpgImmrJH5a+BGubfT2B9EW7aui+3m
I7vRBultPd+h0wd48V27bpwFOd1RG5L6aYzaWW0870fG7DicVi2P/UiJq7NWXHTjIU6RvUo76n+W
nVIOmcxaofADkjC4XnmTJ9j2V11RSsjQOyI/7C6dyX+m6COnL4xQrespW+qWWIXbLKmyddVT1B9E
lmufrmorjPuBts0QJJ9XGi5iX7BNMP/uYrPljt3X9rBQ/PYj46mDyiNmqKBKmkKrZmsenHCgNsvU
REarzYCTOSHRBGfVGI4xfXhw/DbSxqMEtk16TJAcQt5pZOVb0ZXef/wcDkKzjrqBdgRNGr5hF6Oq
B50T7oR7uIv1O5uhaR2Tjjc2iPovfUgoH+CZOq44Xcx+N1kEXELUmATRdQVF1WyrSrN8uNjBuvm/
7Yh0M+BpJYJCLZmd+gN3YXOgtpncBuEwL8lRXwrIT9mortpLvCVy4Vv04hHpacVI0mXc1KJF9ox/
3dDccfwCvO+HqwwKeC5gEJhNRkezT3OrwgCEE9qcmRFbVqvZseKBEK9+mQ2hAmPzXjRGLLKf+Vho
THsLhNhYrnZx9/u6UoAAR+wQepuiTOdSVO4IqbqXItmqilQe8l8XUPuJqBm6dwtIXBft3nU9cE88
TpDqxEcpouQboROdIsOPgv5YaWOX1/QOc5uhCOUNa7wja2aqfGPfdpCPl9sn+CjMZZCOyLMCjQ9g
xyBJa1T3NJ6c4myDC8d06sfufD/cu0Q8wx6UqfLjTHpDpK1RTbI5cpZsdw0NbT0ejLxHN7+FMCD1
RjGcAMhKEN/CZIRCMm6mGmv7zIlHaepcIuQ1szWi5fhZEyc+rdOo5XW5fR7OgA4ea6MYf+iWw5k6
C674Sje43amdwjWBCXaQ/k6C/ItaRDoQcPQ7ZbvslT5dyC0LALCVzpmXP9HSvmbdc+xrSoE3syU+
rsUKDsBrtsgTBagOTU5aHLIXKOBoYtUVAfG+33IxLqBVsa9kpUUPWVgcTGcLPPvA1pQgjcA6O+si
uvKnpJu/g5cjsdV+ibr6LG+BnRfDZPYTPbyn20IiuwjgBRF6KqwxJX5FfGILB06NpeI/QKjH9khU
Dl6tP0HuEPTdwiSRf+7TI+3m8ns6H42fTnLgMvOfwusC1ELSxFeohBrNTN7vhqVKKbYto5HPBGLG
nY4PhEXb/xJlS6aN7UPWcgpbh0LuLVmXtrUYhFuxQAuWr/zoiFT6sB7adKtctq25EDM/YY4Bw0Lu
Ii7VWcIir8pN78ox8Y2uT+qB6SqFHMsZLs3pgIA3j2fzfcoBD7HDo31TvgVDeJTI9q3r6FeGY74z
Np9OUw1agsynyl4mx4wdxeVvbbWbsxW7UdFzMGVKjRKX+gYN7RMfgKPbhIu8N6KK7EZ21jPpv7jQ
pn1sbuxXFdK2+mH/406cZ+IYlGmXD3JlZAnO481D+JskMtzY+0NLX75GTTpDTsv1cqMlLyuNm27a
E+n+MN3jdb/wso2d0BmBVmEIa0lFunDW2cEUYXrreW2W8e3EqpAs9j5kRAuyU5MyTag6RQQkPjLF
Zcu2Ijryrv2GULNBXtlAXGJ614Mx8w02U23EPF4Esc3SH9aHK7+9goD05XbQdYG/9MjbrKIpnp1B
TPqM54dmtisXPjK/X9GFmxVIiJeFi7U90aQzQ5X3ciFR8GL+VlAfvocETxJMdASlkRorYzLgmR2G
YiAbcnZfAlTJ5z7BjprmU3U6Kt5kelrz7peSt8KZUZ7sxafzDHB7pq51H50YRpRc9LswlzRcAnnG
26mmNN55FRhRsek7X52x/zBcJaSU7mSTQOBeyj89BdnhbyXhwwFoay47+xe5oqGu9OVxuy9UWvie
Ddrx31S1RzcImNc7bUTS5Mu4osA07vJ/SJCgWGTxLRf7CSbrJBwV+z0XLFqnSMXM85160IqzNWAF
lVW1stGCvxbWMnvfFsuI7fsqn2NJ0r8NvcISlRcgqWw2QPXg33/j/sIUduM1jv55Xv42WL3nY66a
6MKj33iymm95umcLC6OM4u8ApWIZjFrm9gHvm+wfZVrBaMbXSMitBGkSFpT0fh+c7YZDSyCOVEoP
e4SDTvWapRiXlmJo2m1dU2QT0WacwaOGR4LUknI6SsZkhqG0NTD5OFskyhxHCkWUbxtzjvcP6eSs
ui49l0rESMa1GhrUxMg3t1XQHT1ftELoHBKs1xoz2vimC0Pg155075T8iM2D2PxrSQyp64jjCMBg
FRp22wi24gsFanzYylJFq34yPzb7Nv24tAjqdv/M+8ZDGfOj/6GG6WfTh8/F8k8ngs847nccQzCu
bKtTOI6OxOV8tZ4l9Grgm5llZ0uiOwFG4J1iR1TLXQDfyG/m516vtjmNInTa51cDyHkTf5zTJECN
cFgwZm0wC66pksZ9TTKzKdvZp5ZiSYEI0zG4o8azWYP1PPEhjiaA/aLXFEemIqmKPoE5Ma1bBtxA
oS5o9gSvoklYL8ufQreXGRzaEkfK0e+V/Ep/fj/4/8QF/DdPzRdZXLTRttSosv4LVHNojtnIK0Ng
y3yEPEn/xdOBBWcS0qaSIygxpBlG5NdKbwg8eyuJ3SEO/96jCSFhAniSmfRcGusSdmgMLkcYdxzH
j9WvJIG0pHAMuyBpH0Fkk94wnoM6v0d8CITOR3DDW8dVlLfD5FI7wjx4i993ctFmMhH9z+R/xduY
OBqt4x6Tz6ckcf1vG0gbKLwYcZGF57xzlE9E6UZT42Cm9U4VImdzACPdMdp9+5Qso4dL9Gpyjad+
mPZiX2+XU9ZmCGnAYX2xkILgUKWmbzOIotlSqLjSFVxqJAyXPLGdDVUYkfeQXp7EtAosUe3Qj1NT
LPTjLdCicI46bcZoyl9alBrNlVjGUPjEqICAoNO2MsAuuYaOFZO59BdUCqdnNA/VsjU6URuXO26/
hBdEE+s2BKKy2Y9PiV1JnonP6JFR5Tq29PtGoWToq/lNLP7ZKqY+ScP58N/bscY68vbL4C95003l
lZxyBQC1/sGSP44PrfLZ4AXP7NWCX24KAEVNjxE5pxHXFuuBU+SJi+Jb3jR+upMwiSoyrGG7lMwK
I2zJMA0dDQ9jk+i/D8JPA1T6J2wM+Wq9EBopcvnV/Tg8ax1ymHFOpyfDMHNAJDaMtuY8I27BvDdU
/rZD0F3af2mwtPlz3l9p9jYwZtpMJswsFXIN4EBPWOKXgqjyS0sEFjGnJ7XpgUBiAPTYEXWzF0cM
ZsHfRiHz+XwCK/duKNFKMN+q+6GrGnNlt/Ci1Wnh+6U5UTI0eGfpe1Px5YzxNMNwyOBjjCgS0Yy5
qU6n3t2C+/a2Fcbp8J5ViFzkWKw27XTgoREf69r/IqSDw0yX30SN6YKKeUL6/RY3+PEjr09PKatq
nW4F8p1ArXNutb+kCfyQ/YFJu6qux4buP191ji+9a6gnfnDm7ASeiqA/TghTzbSUUHYLh2CQ2ZaF
tnHUbz8czqmmKB6R1LBxwvMbNiTRg47WkPwbNwCucnQ3h8dfIEK+soblNRDmZGg1w0/0jYQRkxLy
WQKxkd48kixv/J+bPmP+ac7XKrCZRIfZpymTYh0yxv04MphayRQpJtOqEVElR1hyW7w1+cO23NrG
HUt3zOOF63rpxutU5azRgDd0K1/2TXPqpF7Ck1q8AnvdXtFTSg6gAxumGdWDzQN9E1Y0O0qdTASm
mytLmK0vPkK4av1KaWriU1wNnRwOKLt3+Yb/uFFe1kfIDPpV2Ra10GOwhggBLl/IrGlKWzpj22/I
prskqv6wVSvopjkTmUFJKu5LAVTV+59ojpSPltynOgS9338WgQ7WyNEtpI3qfW91gIO9rgZ1DFS9
YJ26+5+q1VUAqb21jnCCLrFbht2hXVFtp+EKI6BR4kQBEGpfr4alj6kpdy+pAt/Ap5NJfIHK+A17
1YBaUqs9WYrhrcvNc+Jo4G2F+fI3z6k3DpyJeGyLW3g1EY9rwjQ/Ws3gk0SGiOkKrfI1le3nuC77
NM0QvY/3xiZla66tLfWH2N2pWQTB8QbwrkWV35wJIb2xh7r5Yg52DUU3JBhzEWq3q3coYRam5PGp
shidanuQ6m9fI/6w6HCQt1zQUANXcN/4FTP7jbSiM5t+yXSPEV0pEgiPfTi+/QDurl5lS8GP1+IJ
KcJyid+3HqkzdPMcuLkbTX/wi8kGXCDWs7b1pokYpgWGjPv6LCBeQVWirBv2lzJ+/DydXWVn33TW
8L7X+nl//wokBRJWt8bdu90uj7apOjlDtM9uhjPmvViFz2ACN/uxlqxKNiZroiMIaXpegw4UfQXV
R8eSijTuJeonp18jE26cJRkJY1h7C8p3B+DVLtj3HXrwo/G8UgB1wwc8g3xvNzdNpRWTHYoeZ4CD
Gip4Yp4iZ5zGxu2Xzq+iPQoxtIkl5bNvPedOo3hPf5hMMn+Yv4SUEd1ztHRY+XkEpxA+Wll0kXtc
6agEhRb9BtBIRZFWMd3wsV8xkCIPQxxjkp1NxtFUWYyegMHmcBZcEOXDWHsD/GqQK6iSp4d1UW8L
QSaib0l+npZkTVuHR4nVn2MJVZkzUyamzreMQvSc6LQ6slWZoJi4BbeFtwAW9QwW9zbpKVZxtRox
Dumm+EFeuzq0ejwz3RXXqefCRck9ohf5CFUrkdzpVN3yR2CHKcwBg09N8bHLorKy255pwITc03H6
zKioBW2Cw6L5FGR1mXRAsqw98Ngna9GZ2qIA5eFs97wLIZNMgiZaeinUhvs9AdbmoibnSZbOX17o
rUuMCUSoVd3XXvWAd7I3G5MowbEj6ATxFHV5HKuxG55D0vDeB49lgvWBrx2BrqpYeA/HStPSkDmv
XsLvrR+tWGx87wXhznWYF5ZgZwbira/JWWDjwSOZmdWKTKwu39r5QicnhUob8pku03dH/LWdLKNe
dT2mqn9BwYTdwr7SUHRvBt2XnOSiyIzCMQgy6A48GYPFQTTrcQ2O9xsO9+SdU3rKZ/Mvxj0OWxHC
7C2hwhJeePJfi63HXjAWuX4loxUqgqWNyc6FcQ+KHKSp55Lsdbb0LKAuVVSlheSF2BAXKQ6Gpzil
l1D0Me3LcyLn7V27ucjeEHBHcq8AtcaxxczY9jFsWeAElEEA42N0uttuxwM4RJgSk99CzeYcmtJt
0vZ7uhXRA7++Gq9IcnJ8qqIw6ZrUHYwVPAwHkRYmXoX2jGcNOvTOyOzNigNERSZUUE2pQa3cxEU+
kXgyc6XWcZ7ABB1HZqj9FWU/h0C1htxhNFR2rbC6hxVH5ivNGFFMFSCF7Nb23VuQhNgmsx7ARaar
bjWNlVQt0YlKrM/5bCulWzcRFv2ra6qyZXtKmAJ7GiMHsvPTZr0IY7x1GWkNmhil2M9h5wS/dtVY
xJtaIS9lbgsKHMMvWo1KI2wk9vvgGb892jHDKEGH/d69BG8lAqWglKDP1cK4EtHq/D3zOZT46sHA
hR0gvMpbVWfLYaqpaQWZX3CDUmCD6JbNCtoBn7gdkEyqXeGOOtIELxG9wiDo9EvYGzdPe/A7rQBN
lbMkagqRAWyUIcxB5zxAAJt86n/S9KeXW+BibnTDAv9cUpeCvWj3kWqDULlSXB+PD5ldTo4AzbVv
R0YwVtgWAtaY95Ujt2P3aNXa4QM0mXs/rq+2o/X9mPo3zZZ5PzhRZvkhMTusLWpIjqulmC/mWIDs
Z7hT4d91ov1z5CS/XxmS0fC3LsM5V5Qx8eLkjt7FbdS0cJCszwGLMLKUWABJvffE26PDYLiFkNk0
7oQS5Q1Uh/3ce22beXOd1JC5yEwmfz1SUiq5v/dA6ZDcVjx3wjbyeT5G0A3rZ255IrAIXH38y7tT
lCRyYCsrC5g91IPMi0uz0S7HbIEejpNu8O7wpERovbmeLtfNmHXWmzc9v0ayvLdVv+xhxxlLRIab
bMvJNp7VAErttNoZ8oteW9ZNhBjiMNQZWtDQNxnIol6WrzHpcwHfLrmuhX8sna6k9c28BdZd3/bA
24rjytn2+0LvW54i6BiPS6LJ1WPZ2qq8FlX7lC9Yg/Ih2029ke1eWLxMx17Pi/B5ws9Dg1Qjs4we
67HtRuV1SjqPFYscqehnVXoOdN9ZwJYxqqf7QnH9swSWWlg9mEicrRRdInMNxhhTSTkSGqU0rLGe
nqt7d5HhrYhiQL04ctxdMjSO7SKoswyL8Z/s1MjJFZ/rGKrMvA7IkNB46EXhGMAZjiJwR83omWrH
ahZVF65PSDgxrQOJtOq5/RZuIH38qizeuK+neE9iu0dJ/5XP4NdeKarWck5EOlKh9jaKvwXsBInB
EB4M6U4CB4Jp1AOqyER3oznq+NcKmtYLIZHs5zHA/nwcQ36VP8zL2RiiJo37L/iDWYoiXHJn8FAg
RqeP5hik+FbNNUobDMDwSUEodfBbL2oibN0R7Tt5FzKfDZ8p6FKMu/nFUrEwFf8jc9NezJFwsj6s
2nm0I0X1LhRo421AIQix0sMaJ0Gpzda8BXpkQrPuPMNFARNpb4JMA868UEdRQiePirRoUuHOZTS/
WmHo9bJJKFWD4HyqBveby0rQmUPO7EjtwRrbwnlDtVdOG1yVcazDqCKbUHnmz3HXTxIgY3Dx3yCj
FVW/jpAQUO//wB+VXztb+yeAC/TLVvDgPas6Di/b1f9TpvWayPLDCEMkMwmDj8vv07YrLBnOeWst
5wA4xvrVVr41ismm0K1IGHm1j52jcxvD/JIWKe6FQSjfLgCzR8bL4TTW9Cj5pD6L+5pcnFrLEg3U
Cf80kX0PcJIUUNvG6ktdN/LYR1Pf+06wztUVfPUFzFcdFevVPdNKaQVao8sp2lLmP4vu4IPiHTYD
Be+7VaH3ex5BSKNnRmOchCl/aBhG8ZzUMxa4tHnSfb+JppXmtAuRbB+rma9tezvWKT1fmMCnnpOj
bCLHSX49Um3ExiVQvtZtHqMKU6Sm/1oRWnEGHser2vOskZX6yHz7grH49Gv1knS63lRHZJuOtvJr
Gc+1hQU0o3reD0hKuAL1QEfVLJpjgt3ekmRfY+UCejAvXnMI8cpjJqIK52XEG3JpyPATZzxzZWO6
61sIpV+XsOAaCmebJ1m7gjrqH4Gl6N59k8VQZjAhCPsoGZJdmpXwPCRLnn9hXcGR4EqJSHfMG74V
ixlWJoqhLKwyQMegX7+IRdwTVEGV1aaSjG8Exye8LxMjkbKkPsOOd71wkJrfZKx1au/19BnJeclB
+85jjUcuSm22ci+7XL+0dNNkLYA5qBW42CBjzcX2JeWMTUe945qMXF5Mk1XadRilRrMMSOhtId2P
P/MtB0uOaalpRtPtIBI0Hp7ElmvYLzPY9Mfk0StxVTrjW5f3xOknqAz+H75BHYrnTin52mSg3Vy6
KrQsGUhdNLtLFy5CJ4iLvKUKGFh7KsALC7tKBBLVM1vgueUXv5YObZhvNC5c0XtJkhjLNZbV/aUe
IE5n4IMb9knUi6eDN9rl3cCrXNiH+1wtnQNXEFdEk9Xl2WZtjJ5Tu3uxd8iJsaRSuZEgBC5tl3Pt
tJkEXS07kZKOfau2bawaEV9XVihturteHhKg33f9TSLlhxdrPOEEbKNXJgOGr/9lRVeauZ4G+WaY
G8cyjtinOgiP14EhpltDOW4HSI8iFe+AG2QOqbOzWg663TdMacUUQ1RXd5RukGMF8F1mHzgwG3Hz
1ri6MxJSV7mgG8wt7jM1lhoKX0GSX465RllgIZdIZELqU2C8HIgoLvB1C2DzMQNpg3WlD25jSPNJ
3QDuIzgFwHz9I484C1ej7Q9V7YfmUuiqu16HWOUWl7RWckqKg7fKKA1NLdLLTcurAqDLf4yY3UK0
sn2dnfNt7jH84HxfnwATsrXTZKh7yaTG94awXBsAhPoGU/0a/NqCCM/Q+Qf2RTd/koM/AyiIE49m
DmAP9FL+HQR4yXrYLp+mYkyxO8P+PWfwXebUFgHPkmO8HgpliurSBeKZZJ4QvZRMVpCzgC8MzE06
pVSTx5tNW7erpSJ9fiYGrCri35abf5he90aKGWdqtp9J31H4oLtfk0Me+DnMBPC5rAOSyK5//3tl
Rc3+03PwAug/IcT1VdbRNqdjDhiQXxq3MopLUCE9Hts8APh9RgIzT1nGBHICdREZXB1y/EXazXFW
0dh03OGqByPUzlszUMLeHqe7rqqn1eEFUgiQaCcLfwI6n1Cxms3vqe8s9fcRXBDfw/PRWY+DJj20
zpwxBX6LZbnv01ypffSn987nSeZF4HzN3nVQ8LP0icSHlLsohiv9hEJK8Jda/Zb6S2VC/c33T5+g
EtiJqbG7wQ7AljFKWmVmZ9N5qF1mpjFhzSXAZRJOZAaEt6XMqc0UdTFEO9D5vRulwQHqQJjPUyeB
L9+Gfbb3gfy8ueDVtVuhgzPSQgkrmHN5L6+k5qw7vtvH5DpUM558vVRfOdeWO6HHCX2bFfnOlL/h
YCGSpxQ75d63yLx+AHlJMxI9n5Xn2tC8cZuccIc43Z4Q6fsma15KmKJai8+0yhgoafVbn55N2o6Y
OpJFXXlrCTqjULSyIrbI0z9sjOLRhJPaiciH31MMM7MRPLHmvYnXKgC5B8TfmhvB2mclWsoRCeE7
SiHyxmjcdwyz/XPapitNyvXhg62qCtPkMy+5XhpClwDOOIrW9rbGJUcd5FMSEZH4akBidpqep7vw
ezB78mdgkK5kpDTVCaYkEgYXsDDhdzCxJPUu35nlJSOusgKUEwnvuN5kI4PyBYf4EUOEH5nxKcmf
A9rV10nk9Nwz5nLfBXW7EMJETJ0LUWiyXRyEPo6kgs4ocQ4+LQXP6gj/isY9Be1h1Vyf3imlzJYi
6mch+WdfpLIzMJQusNGB8QbfLumS6UcUV9rSC6dE7qGK/zd8KJw5BemDZRmRvWmfBPuQ88Te9o74
3liN+eEz/NQt7pb5wkn0uzzXMOoFnhCLVEBUO7h8mqNOdKrvEIOBr7xFIDgpTdlQXlG/d5ik4GoK
bTq6R9PcogJMWOtTDqRmm9BU7IoEMUuUymt90QU+yYEevFwS8PNH9SDl1a5j06fpCkRb4XldkonE
PJE8V4R3KeN//t4gzdK5bhl7+9JHNytJ+D5TCEpRMSlNxmDjWUg1uiyvaWJlpLSikuPQIITFyxad
FHjcP77IdymMK0Jt7/oI9UpEUlrsI9Pd9+7GCQM3zTiK6wRyVXzapkSTFbPRZs4l6skDWEZv/PAh
ZulcTLeR6ZbtlmyEBDkymabX7FH6KPld/LZEwoz6ktsmhbOxYvk+rqvfydIDB2W8tItajTy2/JJD
opAXvpy83JArYfXd3miRTWgeYIxIYSqsjwZ5hCpBEDVtszDbF6Wz1f+E4t8JnE/uJdmhI/QdT29Z
qmt0R/x1oPDHDlZBjKN3RXPAWXcF/qoTS9sDr/bZa7UI9ef+ZqBZJS4BufKAzQ5SDQ/ElCfa5cbt
KqX9MJZUHnlJkxyyH6bw7WfAwi6dwaE4UCXyPDZhIzBRX1Jx/yvum1c4rFBGPJhQ0Ux46PCCuEKZ
sLG8f30/69kdTEdba7OL4Lasvm05DzllhfgwcvMTE7etZ+iaf00bnlm53U4JJXmaULSbRqkxdQq+
XQo4ha1MrYtA11qmKLyBe7P4Nj9oo4PYOhgtFaS5KHiCWdL5CZIBc6EOtZl0tW14NVnX3z4+GqHD
fptAa619Hu7arb+StHKQMPh27GZy2+n49hYTQBGv1Ky6A5H0dXfmzRI9z2UG1udc+udZZwziCqJL
RV3CdlBjszli/Tmote96Z6SjE/8sdAmcdtVMSAWqyqmY9IJZ8GLqSZl0x4f7q1UursSaXMFreiIk
zt33Q450rFWR4pefQOeq2q+I2xQ5qkwKgJX+exCuGu5NWQ/dxJ/gox9g5g+xjflS+v3KIJpoc1nb
vDbs/2b7fNtKWv0gehO/Q1M9WJQij6+BrpfiDlF6iIhXw7770B6nmIkFfrpAdL94rzcH9TDA3Bn4
R0wBr2q3btd3hix6Gpc8NNdVKwU7NyRFyNt9nSslrw8JRPoNusJ/lyq2NJA/uBbvbTKC0/NVzEy5
fumCyuUY8DbP+n0JMVnOt20hdqqv7XbMXm+GL1Z/DRkjKpVe3Fur9U9yzuIkPBdureSet9nW+UTC
ovxciA7y4GBbpW/M1D+hrXLXMrZgYNw7wNcB22YVa39wmr4XdYNOexK7DGv6SzYmT9DnlKHS76Cg
uJA2wKPsobRgTsR3V/F45XsKuXdlzB0WC3tQzT46Ye9o4NHBMcpjYmlR4Hn94OGaYhqOi3x8aNqj
cF4r5g14+7kbEQRg86Dnkrx3D44tTTbAf52Yv9e7GUscW+XRQuOUy01sL844BITgS35rb40F4+iq
tMfwWAE/emOvoZqiBNWrncI+/HdrzB7pSAJNeUyrABdK6D+FYppcPc5jhe2zPao1yix4abNiFKRJ
kmKNd6zmz5SWFK9czLtaAYFO4l+PSiStHwcW/+U6Uz0zf1+i66ZKkBZ96SHutqsBqhReHBPVl1LR
UeDAGZHutgNI83HKJRb9CUzoHFcbmFNzjQK4fvWenAfOL5YE6CmrHl9IZ67Is3m+c/VgnefhGypJ
aHKyyELvciT8ecXM2gEylWv/e+ariwM7vTo4YpmAOT1rm6bMNIz+2wZeR/XsxhXDsptGEZmkeBhR
W3RFV9z5iLg8q30eOPn8fnniCycjC1gqrG7uliz7/0xB4c7bthgL0BOWRQY5FPstceY+hKm+UDrM
yyq0e2UOxUxmrqlnxwt0o4IIuJGBmu4LghTqxx9XyY/PAg9/YjgCeRL33mDErm9h9CtJrSi70wNc
XTBvqeOoWEwf0ZZ5Z4ogX0HHP3oY1HoxBFDSLO70a41qq01w0xtnuFSL4i+2ul5mJngzr2NOxdLP
qvoE1wB/K1l0DHEmzQVtbijohIbubap0updPaOkd859jvseyOOfL9CgOSWj+j2P0jZbAJIu8CdQ0
Kq9mYTglW7mwo7ZJJOTlTko0cQ5BbBrbDxePmXqwGdY8VCT9ReYY8dcvqSvOwRO0Bd5sXEb+uTe8
1+f99pqDfdk02CBOmij3VwkCvCYUwI2AMFzsUeSl+dNn+dl7C7bvRnqvIm4/sKC2h4YXDVB+eFH/
Fu3GCvrMexkn9QMngUdMcyxQiNm/82KZOvODcJzjiHFUXSyMfUXT00e+Ry2KxmJ+Xa5Ws1eBo4Oz
+Z/Ft8AC6Nm9TNhsca3p7dwZpf+JkQ6Dspux/dQyBPHuFnubaqvknreJ++gRQYnRnatJ2mNHIO53
gc0OI9yWo2Ybfq+SP+kH+KpND9VMdo3BPRjKbKP4sFX+8wlMHWRieg3B9rlgunX0LHB3d8tvOoo4
FtUHntgqZU/VXglGnts/cherWCwTTOoJP2KqP0j70Qr5cq0GkM87vIjz/u+079oShJFoWevxRhUU
B/08Fxq8AKdz7sn5dbTre8VGK6L9gzJzcvBKjn6y8MNL64JbDXVzCWjYa8md44Q9L7/ATvOsT0TZ
pgr/6uUlD51AvKS9iYYjbFhc7F+SQRoJM4vytMhY/Gk0BiEw2KrM12S14YTMuBx0kRuvTh0khb3a
Og6oqbSsjz2oJjLhn/UYGEN8tVGh2tWdxZgBEq8lv8uhQhm4QOKCFBdD65wFfiy3Q3leuLeKqD7U
daNcbxWgW3ggIcneiSIfM88W0Sj6QO+ft9QZSn5Q9fmRoa9L9yftlZT19588FgP2fLXUdB4nq6ah
p0bNJfbJE7z/gdji+eGNXW2Jvc/YGa5bm8/jPLp7dMluRVtC9PU8CHTwVy4ltajoxNcch+mY11kr
ZU52P+S9uvVYvdyHZbk+tjKxw2YXGNtMakZ8MP9rVHimmAE8bUkSUa1O6ZNMHeqR+Q/4ernD4wVV
0rBoHUlZsZRd3lQjxBaFPfMyIwn6akbkuyLQfFduAMo/0VRIp02NWr8XnrcX6T98CQTlOyBMmAUI
NFfL5UsziNeZo0OZr8rHugGjkX2rwY15fVNv5WQ7jgVj9FWdP1m9qOmKmQdXGLTwb14IldNgzCYq
1URP2Tgz3cqdJbSrnja3O6nAP3ftyYqIy+TglVFKyoBykktVYSUUKiHAKdCP13iIC8ZexzwrnZkH
gXSInGHmVRrVMGqRaliQVOyA6wD56kmWSqAqiS5CvVq1+NP+/kd0WrY8u3AfEHZDnJ1NNYs+AYqb
BaZYU7ASnKBTSCho9xJVwnZ9chlVZB3JasgtB5lFe7/Hy8xZVEVJiRVx3SksVr4r4mrkdgoK39L0
d/AXZmnmm+wecQ4xg4fOT1ntYyF7C7m6GKvGS2gytxc5+5RsyvvUfh5tyLCQ8JQGMMbfCbEO2JSV
kp3Y340mX368ytAgTwBexFfcwYU3U1asZAdhSRQJxvIPN7TgSSNrkpwNAbACWNv96FLwaROFWVat
EmenCKko61xuUcPoNOf7gd33zUlGB1o6HmC+f2c7+DG0KVf60/7nS9fifVhUCOlMGqA8C9sOcLVY
uU8V8Uq79fKXudbLrf/zGja9RifJxNkI5RoLWKRHKUAqVPlIx60eTx/dpuNXvTF3vWS49uYsUTEm
ADCtjj3NtciAAOIp8KPjU33dYjUucZWuWMW+IGBE23SNarfxEUFlAdz47x2ZAX7/Nv8Y0CHUmXDG
VfySnpbLSQ/5F3QVcdaPlL1KNKVMSyzqx8lyCD8GoHT4eriiZSh+q6u/lmBXd/r+q8SyiiZl3jg+
EX7NRXYsOHk/9KehICR6RetCcQtWPGuTnEunYX+ghSs65CgO9CfuXf+SRuGw0mfh7a5hJvbbOkRo
CK3C1u2siph4RvLMreWBsoXtZPA0PGGwsDoGMFUFHtOiiceQCaPy/5XWhpCRj0z6y2jL+Td+FAwt
V3H6ThKrSIaPUZVz2q1ndaZUzmEixxhrlQKI7tv6re52Mc+IWf41ntjTMajotJTI5EVbhsOUG60a
5+KD9OMY57l0t/Gdwq44NEshgyx2IQ0FsSHhV05y+UIwgji1sRpRuc8lzzYx+DkqB2A8s5TvZhYq
kmlcuNbFZk54IAi+hPojaXksXiNOe3/f5gNE+HWFdKTk6ko65eujQ8wdDqFPj5APleDvIrkK31C/
cUF/hZw4GAqH9E9zVGQf+ETtDeA/HoC8c54Y0GKo33sAMKB4NzdgD84saqy0jkm32GOcMnBXQNS1
5wF/vLmlfsLyt9rWPNSMFl/QpFq86yU/KWETGma1WUeAL+6q7lO2LLK5jkkv5KNlwkvmIMaZ9a/8
iOMzPYWzUrWpAz97uaRGR74A1fIJhkTsre45FW17DX7SUQkEDg/XaWn9b0du/eVOc/MTWrQGV/7V
G2bfJ7VX/FY690B+0LkDfhTj16jtG2C3NBwYIRxSroYhVIe7f99nf4iHM1wPY1rraKDqIHwhrn3L
+wFqf5EHHAPKIXFbiWFKkrEluvDmZKRNDVbyQn7qQxg4FBmVkfN0oTxP4cXlYhqTKEXPstpfgyMs
H3sFt/+3Nm/rczYpZaYK1eltUp79q34XX5HR7xxPMwwdUpr1foH9HYMNhSHLgGKXl7qVxqPwkPGX
5ITpNhGQ1YfkLECQKVDPazfJlDhbYVgbzm31w4I5AZx254kvVAilmpKyXBlapZaihHnFk6edEg+5
Q6vD7nZv+hXOpiWEg9wfA8y0fXar/iVWfGLqKObxgmBn9BHV2xntZjc8RjLm3zqQv8N6CQ9bN9ht
2fvRLIUs/01pwPS600gH6gXcTHYk7eI+PaCHJGk+Dx82vip6vPqclg7JDlbpSGnCinEw+oe9uy7v
2ABMPp18ERhT+2qgNftjQ2UO8YxJr8C4etQluIYSvP7JDFiiQtf+eTvNYPAD4SGniuBYWle6luI8
c5w7ryNy2yuY8qEGzcLHeZYmPlBax22zocQRxuVjnIL37Zh43ZxZSLy3LLQSt+WsVUH/smdatOhV
iVrYYIBNteaXqvziykE/qHYedAuvOdhz4PHBfC6gTci4/WnBiMtySCj5QwA/eYv3Bxb5Svm8t4LE
OY5llj6N6wwOkY2PmNPVli+GyBHM3H8MDbyeso2/NM0J/ndro8fZvf+rDTCer7gap0fUcmQac4gY
NNfJj0ZnKjhceoVCkXAubq7lPOy1URmKqGHrZyawyNXnT1zBGcKkQACrqKQOTgziT7RJrdTWxKic
D0QoKwyM0hNrXQDC2lOGdo1lR2fp7iN5M1swnU678z2U10abykQTWNKwKFbWJDMgZbf0GCYbnBrd
e4MsjLm8QHwqelzxf8RzyuOaaUbFNRrbb7q9OxRLXcm5URuckkARcBYINWMviE8Dyi6GptBOassE
UeezeJPVdJZ++u1ZP9qwJGmJ68CXQ0SxDNw3J9mAkHBpLaui43dfnT7KwqPq1bwpIHkj8RI8RC3h
1DWU1FuRw+0oK6h42J4hML20qXzDdaCLoOp8gSDxgrAxuoySnIlYoECUCzmuGkfepXIuffr3spt7
JM1I13Nem3IyV69xwI2KSuz/H1H8I4S2O5yS82EbV9R88zA8oR3rmA9YsL7IOh1RUY+/9J3Nz19H
DKz7T/GMwYfL5RBesKIf2QIB3pGf0cGO4q1je56lkBY49WT5LPEyr4RRMxHnXEDRTQUCPIY3EHi8
cF7EmB9R8GundJ+Zm6GaFFJHPqRce9ObyphypIysJRsc1EsBDfqjWFOoSJJ59MyP66VZQXmmdoPk
LXD23yRXZNKpV8j4hgEGu5dUuEhp7T7/cqVhSMIKbCiLQ1ebcSXcn0aF6U3RhVlK/iB2NyrpJJW/
VTNnPoykHUbIvHDCLr35XdW8luB13/biGRonKQPkyGj0UkU/9iNZd0/nQNEP7wJtCrAyuV1nKr51
077F3AjtAnFeZbwWzyb7zVW6KVeWrbDQniBrH1GQlDgklPfdMH9JCDBkHyqHaDrVSUhwAZ7RwliG
h6jI69+maDo3Gyf6pcfIobtvvouwrZhLyIDh/Ie6DXUXXRGLMiK7D62X/cMkxfTArOjvjonmlbKr
qAr57GLBuB2BmUQAayvnJt1GShaf867P2qpIdvTlLwzasv/IEnHq8bKUFlvJDkxCiuRGHgLXkeRv
1XQLLjs+PIKO1vbPQN0Y5BYORY7PY8qoz/RHAqOWegRx4kggtQDnIqZbqA31J1gzelfuVFQGxUh0
N6KyZe8bssBX+g2Dvm43GNsWeCtkt/6P83i3lLunbJmS9fdqN3drqD/RGItCFpIkCKzTveK2pfgc
fuTWpRkTgYBUis6DVvw8ZEOuAAi7DAeOWBAm89sPOslygIBAa4NkJ8hz44i0StrEp0BockJiBStt
e1TMZi7sNIIDudVnSZb1Oo5fmlboZ6XkUUhXop5oKEKB9umfMPceROxjUqz3UUhfIF8S37CNWe96
K/r8UwnROUgmqtKR0viGgR2kloRN210/lZCHpLRWVwRUhzAgqIz573SexTRLxCzievLp1Rg9A9xL
zdqs+gL5freuZETt2MDkzZWV19wDDQKCMeUXhcUCL+CjRDWbPceaAJWJvBh3/UVjoH8Bxj1nxgLz
Sl8oJsM8ZHbYvPJ8TlRzcRFg2BcDWomKCjLXbD7ccRVDuqJedDEpfTY6vzy6kaopbOBjPd2YOZc2
HnYof6uXbihqEKoL6uziMlx9VS3snpjfgFM96Aqf7zH/L7lMThSi2XtdzTzRijGrXe99sz2lgNL7
gkej9J/crHhtFvdubX6QFWi7h8CvU//pXsp7+29nUGBQy0rdf7VOf2GNAaN372qGHc48Sm91SA73
9sivxeOx6Tm+wvEbdunc/GyudT5Xk9BX7Gb/rLQ6zjm3uF8luCp9x0axn2joz0D1teCazneh3Ttm
rbJ9rjPMgqH6iV4C/3985Qayc4JAfT+N6NavDsrrTZEljGUv3/SYoyu1jRH0It3rDhbdr80mv3pi
vW0JxvJtrWdpzFAUElu9BAQLCPbIDObmGMkocQGBQkAS2tHCinUL+QrxBSTL+OZQUwuUjPxYfMnL
haobDljHZZhxatHcxtz8xyQ5/x9E4mZw8OSFNXqI+xDrujoO8A6oHehEYZPOb25siJzS57nUJYNL
cEaX8cKbAaRTKIte1HMdX7cKzgAhKJe6z+etEXtY1dM9mNfFMDB/4lJ0E9l32CQuOghZnZ3ul0Fe
X24Z9p/OJMSR2AyMO1Te5XWB2oNTWGr/mGYxEtbkP7KGvPBhOJUdCJjWOZSaJkd4ENFAXXAx8VmZ
pufQKrefdGBcTyrSVOWeOgRFY80U4Riar1ZwtktC7JPkERItW3VyRt57gR/YEs2ymKiL8EmcsB3l
hD9gWntIXoibWVQvWLxy6Qy0PlthV701/KFyMDx3NxHPM2vFX+FcQXwaZXvcZby2pHbnrK45U76t
67Pi5T9TgZclv5WTJvs/ZZwUqgejTdEWaxhjPehNqm11tt2BAbtBy+Z4q4O/EUHchF5oaBfW023q
DrsAtqhq7jdmoKZzjWVo8xrzL52Qg/ViECTzGJVp9AwGjZfcJRzU3bwgQLDyqXF4yX4k85l5VFdE
/18aE6vt8ZUgfm40wUohnXzBLT9+lr+BASK0oKupdGo7Fid1HeqaomhQrCnDchJ+v8aO5hN1mViJ
R9LSJKN7Pp9PotskHGNFxbr8Kw9Raskb407MgCaQZGZ6avlVxHoyAJrPyGVbsyXxWfcI/ufqtsqm
UovdEz4h3rkquR4EANkWcjzkJGDL7H/OQHm6zQwIqMT/8eP4vQxMG01tda3R8uMf46DLufLuV/b5
0EC7AIrw3JMicnwwT3CrctCDwyfaK/PQ/zQdrzXJz19n8QLcUi5PzLaqc1t6QHMQxxePlDnVAY2L
XqF94ZGnddn5YpRVo0Dp9xLo0AhYI7ADY4HmD6p79JVeV2lXSqwaWfPsgaqelNSw2CJflpAT5nI6
g87FISlt9SpdpIf4tz2Gg7zu1xbqFecg4i335j2WE5iJtZT5So74wTNZRWCYf4vrWLAC3mLNR3pE
mp1hLHMy02agkXX/IfOGtnoHEHuSC9gt1y5ZwEisaPbdBN+tc4Vllc2qJQOykyR0dxtjcBgUVfs3
Ga03yNZ+Wu2m7KRqRVF68yX+iT7cVqhY6LsxsDNpJWZmsrs7CGyJ+xLpjWipubdiX8kRDef81ruO
5A/7OthwlKgIdGcEWcHnPwZfzpLVFaARjDvP/EmbKQcPYkX2oGQaN+l0pYowx4BSnLm6V1BxZHe2
TWN6zdY1xbfN/m2AqSRPDSSrBTtl+AzfaUAfNtRcKub3r8ztxDBZ2JJsBvPwD4kJw0QoeLBeTUrE
fzJ2R0giAOuLd5wKozyNW3+B0hZq/1sY4hA1UEL/xtGsdAtqqi6ocwf4GTa2SUmYR2wE2BvuLyzm
RbTXRnTpmd070ln5X8g717oR9vR2U2aoEmaGyWa73Shp/3DlnacUbWA8iONyZyWo5qNh9fepKsks
A3zAkgvuoWL3rYWMrTsgjojRpqRAMC4iKbs6E3PXlqxDnXLlC5p4RT0uvFkwwB4bQhMoKMGcMNT+
sVatn9w+3alWD9G9lTezFvcGidamS5fNBlN2vApNuY+x6Vdxiis3trJHCPuL3ce+G29dAtMq2tj+
O5wjWchkkt4/VtyBc9dNtTEs9RUKU19LLeK71aNGSaIZlioRhMvcczyRhgbL1J092PWJTdHp59MZ
4FPUv1bYPZnMsZkq3PhyMSHgloAw3QGanrug2CwL0MWSLFQUtBV86uiDsFJmQ2K6kBUIowuDYPcT
Z6+kgfxdjRcdQiVq1+1IQnUDpXWuzrzqW7+/393fstU4dlkEbsVYj4WghUWn4SMJ1dXQKJejygqK
Oo74y8txB868WOXP0MsRuMH2IhDu6GW2GmB62cPIgU3xOrQ87T41ok2/C/fMyxqxe91oHFalORV7
6echKaA8TcCUD8Fb+9JmI9bhtwWGOrLahqMlchHYdRrIr7wKQkn1IdB97i+SguDyJOUrv6wDj4Yv
Ss7C3SDVH3VMj0OOLU3XxxdS+8spP0QZ6ttvK86/x0VBI/0qnV855KAE8S6oaE1jBh0e/8bw73HS
6SpYkuJwDtUz2cDMLEEaKyUCeDRWkIVmLF56TsC6rsOlWvqPLQ8KHX0CjKAQDPwJsTqDSDe+Q20z
MUz4AfJU1kr08TPn2n4XwQ+0mg2sWzJ8s//vYpYJmwuWhsY7CAgsINY35QkihNyAd97MukDH2fDa
IA6a5afN6sNf8uf1KRNRPzp11gW0NcOArH3pFogJCtcZR+3x7rmIKj7Dp7BAMevkX0hbz6IE6RNL
Crh8P5iarhHZ1ZPbNKgt5RuF2HneTFjOyl/H2+Xe+slEe0SCRCybpl/COQPKvl1b2bTbL0n3Cis7
FNvyun104b8UfvXq5w0Tj2HIZGmFHMEt0mlmcbqa4Ofy2lNL7lbA7CwPtRI9r0NmkHXYfw1vwSa1
jYGdl4vhxkpc9xQfn9NUXba6Hse8/eGIc705dQG7yO4gslbTq3sWb3oCHGgWyQ2tDG5HocfAuu50
Dha11osRdOryMPXi3ZJ3K43ca9Cr7Iump1zMfVh7+e10+gwecKfbKtEXgXrRIUDeh8zPmJoFkp1K
44GpBzavo4S+WSjL1P4MuuZjjojoQIkvA1EaLdGvnMYiL7rUKRs9CcVNhRvb6ohpAvjLU3t7nyqF
xyx7cc/VMZg3dySvYOLXPu7c0DcJjUJtguiV55E8Q7wM1WRBUw+Lc3Zu9MT6BPDwo9Dg3rvKDNiR
76CPddajNLlfLwCUdFwJsMTaU3Gf2LWBUoiXELPaLBhDL9njHyG3LKqgegdR29kfqhs7Yj1TrRQg
DcQkZNVb0VX5DLztFp5FEGXTJaWpYj044yKATa3a2A8MRmbrYasK9H4LOjERPT3bXdCbiVriiCXe
au1zbIkN324V7NGADz3fq6Z7g6kPr4zqhRBeGSmLlc3QogTjl9PdtDy3th2qJfcU6Vo2fAghU+50
TEZV9zaq4T8HCuNiBr/z0d4vtns7FGHpbmdvl5rd30lqsHX/GesfrEq9/PQ+O36e0hUrToMeSVrM
7F3lXCjaNvLNLpaVkDbq6oS4LaDOuHrIyMgeD3+MUp5lfnGP4S325E9qz3uL0JTEOjshaP9D3cqR
Qjpvq6YQ7kLv4W1q5d/AiF8PYetzBSU33Ix/0ABEZA2gvMvvrB9LtUJDa3hqMZZTMpdsO7cfkkJC
dfkmq1VOCo2YIE3uouIgRhUPkSN8Vqd8pwNp0BgMnC9okIfGJ55qES7uwtYiAwe7JKJ+XodpTdZ9
DhRToIudY4ywz90UbE/rl2g+StRK6XpeYyacbOJXNtk4+GPdlGuqQqBbj2YhYGV5Ri9KQ5j5YriD
U6eEfjIueMB4oh5NBmmeNlGQewWFgYmVF7ztCSoNupyDvHuIEGbvNMPUk+l/Q+l/zr0l62L3jfGC
e/T2ORMfXm2Fu1sUzPwKzdzuafDUekQYaEzCspyelG8JZvLQFJ+POfJk9GxgQgT7kexmjfbxCfOM
qo3iKbV9w9l6GA4sC3oxguYSoX3f/sMeRpcoLh/MlfNeZJaqNxNMbQ6gEjERB5gWCUc/66iMG5ez
gQU73qidxGMtI2KIKHlsKR+2xIDQyOKhM0ftBQ1Z2RB9Ac3HND050/fjlUE7tvS/I4RNawEo/HzJ
UoOdzB/0mv0Dq0z2CWttmx0UmmCVqfleAF+8iIQtqeqgjPoymkPmsAO3YzcT77bpXq/ReAO8qIIb
AebIYr5xZI34EGYqzoCbBwE8m7vfwVdCtEK9u3bInia5GfWytfbjDJJjPWAX2s9u3wm/3NtzyFHT
PCBtB1OtIINHPJPOaGJ8ojzU3/1VWMkggeAEvTVT7VbA+p7pc10eKBCP/IqD/AZ0+FYNHbbSu13+
24gSNpsOLhOIdeLy5gmZDHkvsyvCeRIsbP3FDh/9TemRBjM6qZ4wrU0aC7OwjveE86nWofgw5dJp
ZxvwthEVifsul/GCpwke5OALpgbp1ySfnPKklwkrcqHgc2A+Rhap1YVqheEfNsOpixarIPWcyxXh
PuVBkUeF4IBgdDBCVrAXyu8Qk7hGGnmOqQh0BW+9o/yyMh/e9nJ4jTzvzTwT9+1dDL+My0fdguMR
33eysIXERRUzZpIRV38r8cyy2twE3Tt6k5ZxTAOJ24l2cvaFmKDzYM7qjVZ03KdyPDA3VXTnwpD0
3ZMkU3cjDzXHF4P4yCHRvBsgNIFuT71evMuTbzEycFWOsZl8MXyDK+Xxp6rJJ7k8QkWcsSt327Kb
OrxzoQ4SDAyPFrfdfk1puupIdhxtHF6PMoz2I+ar8OJV9sx2XJlGL2jIh3Y/NC1VJW1ao78MkqXu
I2dTow39Np5+h8x3efvnAshJoLpLB3xZO6qn67+VvRzw7iMHivwPpEkHaMEqNxkL6owbQKve3cl1
0IyFS93ezkuXiwFkw/zmuln/TzvIe1ma1dPYXbu6NWrqa87736+vHzMXNgIUmjxq4X8Wp1bCqD63
OAvzoF36ttcii6nDKUTw2xzdIuE6qmd+SHlsD30l370GoIIAbSAeeNl9BgJYBk0mo67fgIA2o5Cw
MkBe0Oxh89qgKiO166M8h8WOnNEl2uysX/kegJeFQBcER5R6zRuuyWDZnSB4AFkR5DHA8YzNxvJ6
yQm941PsfB6y0lQkdPj3F/MXaQx+U9UcFV2Q4pDmq+AztVqkxKWY65qiQXAwWMpRW/zdkHM7HnE3
DG/8SDprkdx7uMuTGzAW1L24MvjpDmByOYllw1Q86wErSIU2m9nqWwWfQi9vtmkU6zfyAY75fmhJ
/vOXVY90RAKkClHmSBud/VcHhrWJmv5AQYZjpgEZ8hFHuXBNH5Ttr9gW2hvCDlVS6+DiCsI3Ku2G
VIW0Zr8df2Z58ZsV/vdIRl2dHFxigwiPh4SKnJ3NWAvUkSNbrojG5aaxtdeADaLSTLxAkubEJjIE
Kxl/iIzRWFna1sZgElp5HnFyPi1FmmmWm7QMOEYA4QeLUpPEOv5l2jhUrW78Qy87YYD3AWubCRsS
dMX/h8RdGnjNeaajl+2YA6nyvVh6kab9W4NvWqZSn0mmN+MDPARgQSlO3PnEtuqLhyQg+39gl2nI
OyKXPpctsV3i11JWM+nOEcJUpEhvOZ5Czgud3gLWNRc0oPEcsZgSlOpKlvDAowMPb1CepwVLj0ar
9dDEDN9E9FXbCSFDdMNEfOsot+BffNu/4YC81/hla4oqxh0282iumf55mHjhEPEMgDCvlMX89mvV
Dp0BFyBt1Y+p6Lx9Dq7AiNcav65n6Ec4anzRsMgPjS29drJpvW/1LkDtYxKh958oLIp9KY0BlgrD
Or2kAVcaQHgYSo6LETsM8kqgWtSfR0JuY8XV1WlyqphfhXyhmUv6VjK2p+qJUfMxIj5z33Bv9h54
dKPbVSDqaNCDk4Ij3Clh9DhYzoLGcQACrplXNSArgNcgVZ1sotWuE7C1Ub8srr4wXKYjtYSoelKs
cXxkH6JqzxjAPWsoycPw4RAJt+vE+1JYX8r7jmV7ckY1khQifYzlnNDvC0uJB3Hbfy2+H1kBv87x
g9Sr61sGlKMUMS1bzHEEEfdMoLJD2Gi0Pm2fBqOgKOp1ZbPMfp5aisEsFIFjA7z33hHN0LFz506e
iZqEJQEMYCwMwJXoyG2vACI1dNH7h2sJKPGGWUUvDOCx6srdDOAqWHZjEoSXFCf6S/4Hs7qKEvP1
CtYeCuj+toChericor7rQRGNsflmg9E/MN98tlXAeXT1hVDezUV/5FBtTSn+NMBGue8JnWAvunuP
A7HTZ6smhWoVzysQbaPpUQUQGSORDEmAF2ClWXoTAueuNDj8HGyxS8v8eNHcHZ/hSEtfwD9f2GBl
8yuzXO0erRne2O+g16pCaxk6LsuUn1To9DHTkIU1iLsCFSJKxQwXMOnyae8MhwcNQXbi8K0MuJNi
uyyL9H4ppPcpP0YMYyJ4VfpRzj6530kSsQHa2IU132sA/Rw5Ns2ZfIsb09A2nx8/R00B/sq5NsMD
OAcqjcQIofoa7IPb8UCFTbiMuSJtuYh9Ytk8IBHNBfzRdQqCnNAJ4YY4I2P6+fiyCUgmuB3Pw6+o
4WWkYS+ApLnLX1FPCFvV/Be9VLEsH6J7Hsnhplh6sjFACD7fCXy9rsywERQaUvSodjgXYYP5kNLy
vxjiY6pYgkZdO6gNhUqw5KSH2Di5kHs1IRwf0iKQXvY4WabUKL+ExVu2cOLZ6nVLL0N02EclLJT6
cb+IJpLxJfRbcls70V/ONl/r7Camt2tSs1JxgjpF4ojxcAX0A0yuN8wAALAEs0Rx9Al5v5/qibaQ
+lDhbnpocr3MjmjZwR/oEwBMwDCiGmolsaOW+77GMlRCw/3+G22uBtpWe3Y9f48TRrIKfDdChXVH
Um9CXTSNXCmfaoP2InBLnswG4hqX5eglANodY+fRPgk4iLJsOhvBTFsHb27EKnap7j3ABSYY2YnT
AgMwxc/Pt+VAj/4Q0F3LM8K7YYPoW50yc7tJQ9rG0MnnxNQtYvAw9SFCUyDy8HUuY1Ptkm4bOkwc
n3TTrkDn04Rn1uEvYxp0QA28dmb2Dt/d2mY+vftHe5MDIXSH9oq3wukni6hS3MnHjO8ddbENeED3
1P+fKjhs7GOdy4V3P8tEJOzQ9MrHLSgvQaSRi+l51/6kzzQuMGL/fqh3P9saSR377q7mOig+7BPR
AvC/SjOdJozM7o1gfFxo9jeawiPrVHxzMrHbiraCMzIax1YeU8npMa5DNd4ueSal7WHZKR7Y5+Nc
1ESmsrzhnYgELo0C0ZzAVacvzibL+grVwRdjQIF70yHptOCTb4p+tEGmQusm/6WUlim8kJt8dgiu
m3joG9veNH8lsoOAgNdFM8u3qgG84weej9QQ3VtgszK11ZjaFaPl/SZyVKfc8nqLDFmc962zVief
dKRBDpO6etS7BQ0aNrOPOo/tM2dtUJLJLTu4GpZr4CNfIjOpt6EI+5dUD9oRGBTOvm9gQtM/ibHK
91WlBZTvt3X8XfPhbIeJkAp+lUAW4sRj5WmEOH39aA2MGr6+LzYtaxsHJZBLFZMdpAq/J2phw/2f
VGd8Gs1k1WTsflNZsRQJHJJ6PxyrHIqF0k/wfgATXnQrHlnlRX89yid/Amk4g0I0l0DDGVX1fPtQ
vOLwfoWV58DDbnGEV4Pbh/KRudGCiiEUzU1L/dSpI14WabDRrH4SNPdZQzLnymp4EPdl7gtNwlX+
ZKKKIU9IsCUwUxik8sPoOSNq9QeOVjEWT9De589rKPnMam2WMsPp16/zd/5h9NQnXN5asQ+YOe28
OHsHnWAGDzkuFibzCwkLslUsW+2hyG2NJBLysIg3n0XF3ADvITnpOoU+sSTWKucNgYA1D23sOLaZ
9MJvHm1o+tpahwiMXA4buiZvj8oz5CIy7SG4e2RMUuBzNX3oufR56RgsY6hyviq5/IzqQ6qYrE6x
HHRJOCk4sjrCZvT2kYtLucUtefJjjHnuU8U1lTv/TXaA5QXY9Q1jssmTi6cUBBUBPEQEFUQk9aPm
BXzIGsA17JqhuFy8AvFqux7TP8cQ1Pg7xHkh2nL4Of3r9sfLDA4uyALGyoC9ARG/9KTZ8ABCkIsd
fHH5BMhE7rTr+gx0b4Yw9jvD1lzduomDkAoqYiOAVvohUq7tJjq9HGPq9hQHcyL2sg4zGYYE/nMj
zwyE+q3gDLmputnrkUN9LboS4Gn+1CKSq1D9aHr6LkU5/q3Ie+et/F/ZovQP0Pk9Kp2By2F/MF97
VAkmJFXT539WtRKxys11Bw1iTEWWIG3TeiKDhYc63v6WhJPVRxhgrP5hrC66JakgxvhRG7ftMa9L
33+ZalPyP9y5cVP8QpS5FPdKL6jJ1S+U8CD3QJF47GdLo3ivfk+PyFxSWgMjMEBUkQlk/LhxsKJz
97Ix5a4EAF5RaUAvKtJPfZW5/c+3rkzpWEiJGTbXfONycwgaIQW0z5rxrltWsPpQSdWxXOKodpJs
K2Ss1VJbGaaJwkkUcb2NE5PuslV3sY+lKJZ2SDr4dqEogRwvdsLfjwFBBSQzegOvIAnkd6sGqCtb
pv1KcRnmrhrbcUO9FXWnJw8f42g112aZPugNMaqPuA2QKREFC7Fo76Ui/VXD7kh007RmUzp5lMop
+1vePORTlM2NcaqMpWuc0vVdjkj/N9LVzX/r7Y+9wBFkAtxUvkzW53ypFuX05wvnQPdaayoX4k8K
G06vbOUp8mHKPTEH/SJ7/gNW09YzqNrf0N6rHU298nEHZSpLLr0cc+FlaZcU60khELujMG9lsAtr
npSdgh5T1KZ9luoD4snpc2nx5OEgC0ywcZCxwtpAdS49sHK3/I/O74AGpDA/xkE85U2ca2A5KOSH
XxKND7s429inXErQGHt1oNXUedcwC+xqnpqDNdxCsZgUAhl8RYUEwwQZNbb0+moGZL1w4xnml+5F
JBFwmFP0QxYqCPizNlDCzBNmS/LHGVnPxeIg/TGo0zPD5ANH7k12PyFUNSoapw/3C4vDTzGIDwFZ
W4ssLzil3PYsN+lOy+LwgWuRY1sFImL9BgHaHo7HSQygSNbXJBdAe2kix0qax3jMJHJQ8qJDQsmh
CifrpfQBrc+QYww3OnynSMbH9ia7f2Oa6P7GXinTqmjQi9Gp0w8edxlRarpfXELtNX4kIjuIYj7n
q8cuT9hKKMIenXRZ41W/ZAuVNa7loScwlQrrBEirpE7WNIzcxSMt8HYPK+AM1xyzUbtQzqeN93Ru
R2z2/5yzIlkk+rrsGkICWkwQxXryWZAvIdiNSzzdVPew/nOINX4NKvBNND84fnK+QyyP+TrEwaoM
DRX4NXOImWGlSSGjtSyDZ2GInkLfISdpHOJs+/KISoFNHEcxZFR5h+fzNk3+UZ7TzN6NskjrHO6C
RLp5HfNOCXzjFJoy6QzE4NYJ21DlfstQbv6Feiv4JBSeXaRfYbI/H/AM4/13bwzZOmIu9tPzcTkw
P+I789d7yDQ6ZaMg1aOojpDhA0K7uHNICZAtZZoIcRlflbBjcGYdjMIx3IhZI2/iYXzT8yRR4u/8
SZAc5ZpwaG0983qhgvhl2OugfUnHk4h7PygjRIFzlf8lSOjA14zgt7ikEZlthe+MUzbOTy2yivpv
mWhj3PYtfRoyOWU1xqYB9RoUjGoQt9VHLLcLq0iSTSmdJmWE5NqNuLpooyptTAi7AUkgBh4TiqlF
8clz6igOeoq2HMPprzpC6w7RPSsyoxGXa2oQ9oY2GV5Lg1nhUzh7lRRLnzWdST9hfojzoAX0FqbU
XHe5kkf8QtdWsWMwHxQSk4kUiQELSp7CpzeGeQelvwVso+Xt3hM7Qg1yFkiZrlgF+C1Z9PX2u9X2
Ie70y+7KxZG6mYMfi6IVzXbA4nQOTwxGXgU8yQtSZdiYUHlL2GoJFjSOW4z+Un3ChUEj0fJIOeQj
qma9lDArLJ606EYLE5cl1DzQzklxejtNJikrlm87WBttr9C6xJIEoGIVilwmJwZYkDndHHKHIcna
Gt5/Jfknqm7JpYR2uy7MZ3ucu8OAkjEPDJLuCF2OxrO7kl+YR2lK2bFHl1QxdUIHZ4fh2q1E+ap3
OJA58lFUzHQzpUW8rp21TXzLxY8lTyCqQvjgZ10J58DRNTyNaorr6yLzOwOUD4d8NSjqGY4TSDgE
D0uOOMHL7cmz+fe+5xOndM1UYw16bDCeOkZzW0ERWYunYiG8qbTxkGavheLVmwykiPEKHb4PgeX6
kJKnTDmvSqglMn+JqLPWMcywieFd0VitYSTwbSnQDgJetbyF4j0vS46Vk1nbk+AgEGJZ3Mw8T+Q0
Qxk078KIDJZPadIi9eLK0lfN/WcMHLnLCMZ1pNzX90Oc0LfcrdkFop9pF+RV2PzvcJMfN9tjbU0/
2gXcx26iV1WhlBkLalJm9ItpRXnPLbltGf7EtfRS1OzOXNLcQ0eI4b25wUyiikkQfgPOWwEQMo1z
VdIrZvr427aUEodAXElNf65IjVq6qxrdXA27edrWmFaZflPQNnQbZegkWGWADzFynm9EDSnUHOT2
OdYb7uMndgwceHAZoCtqItW2gKVvp6GjMZrOYlUmoPI6C7ramuC6SFdcVN/ecVpYPaIb5YuA8cx6
6MUPGGfIrngET/saliu+4Zv4cV69OJoWGvnXVfsZC8F1Q0K6mBHqYHOwJjsmMjtrJHKOb7P13Cyk
P2HqTdxpeHKr1bvABSyv8q2pDISOmUennBZaEg3j5fP8eXhhShUwnT7BjXm/GxVtmIfthGxm/U+g
D3HKiaK8Y1HQXotwgLRJ2U52KnZjgJi6qBGhQhWNixHi/HiyYvwnDaONoz7KXptVJsEF4X+Gqnp8
CQMFTN3t0Rz208JGTyU7CIdhivp1EI2RPk4oICFlmLlgR33e6DepY+53K8nXS60/TLSHeMBji/XC
fPA4P4YScXD2/OOYewYRXYkCrqkNECeGGhuWhHwQ+g/o44GiVIqVAIh4BXiORwnKfqEhwr5PLyW6
BK3q7hj/lN09/s7KWuEQPA5YWcBqKISGnaCwMD+O4M2w6jD+NFITAcMTc5lI00VDjKGysDuw8S+4
lsVvG5wkyL0ol4BCftDbsKapNw746q0+j1mQxyCOnCEFX6LV4BD+QJeRBSDE+GIYXXEUU+8SAbcY
PwNYvBSiw1wK7V2p7YwYpXEwDRTEB6O3Sls7vBqQ5f5dSVDQIwo3ggTD6Z6vjEZ07Z+6PZvxP0aG
QZC5SDSUpez5tqSosFF1S00LRlzvkgA0eK+u7CImuXqA0T0I7s4Ofa9jbidAKQpCz1e2yJ/47RnT
JngYqfnoiWuz/AGuZeRyYMWLcBqpXGaTQ2LsnReBdMlEHHaCED+FXxsrE9Xodz0uKLwaS4vgets5
a7pj9hcAAX8HEKXO6msxQwR2SZ65URNBt4xIc4dIx9rJzqgiry4FkNhQ9chDT3YRNJSNeg4PUgce
n2gqrvI3w0El39AwcKgmS5v9vHRXkV9kz9jqnYLjQVP6wcB1Cpg041GT/NX5T7Dxj85JxwLGbMIa
AL1Lersl8723jkEybPtSx2WI5Jx4zJLNrL7Kg/dZ6D99DC/tXwEApkDQw3v6Wl5VSQ7s8hlnLiHN
12/2ZRqxs/vUDslUKH+8ixCHXe5ZOjDDg5ioXuVHMU5O2r+23O9KNmNm0Oc2flAXHjn4nU4X2g33
bdISK4vLP3wWOWharDfhlqm97VDSidb9LkK1GJ+PPuNfID2LExmLHpzsiJSqzFaBTl6kk/TjyIEO
nJV8DHCIXGmhr3ZzFWEojybQsOdkS9TB8pLRtU+xuCFeQlWWFMQnstGPwELbKlTOfrndOXtmW+K7
37sIeQsBN68GatnDXGMOga8rPvZus9uL4pS1NJ/VksCWimmPN1Z9cNYEfhBkcw62/XUgExX+yU7X
whz86ZSTi9GE3ZctKGWNTQeaWl5V9ha1xlYNiPEU5gpoVZS6PN52SensnZfvoPnZWmH+T9fDUgVc
2LNq/sIhJ4qKUpn+XOWEzQXmjLGFeO8mXbnxBiWsnZQdkeIWUYws1SvYwu7xZldqV/FqXpAwHZcJ
wrb7ayrTEblJEsiaDVf6oeoDROYDVgO+EOW6ZfbLwxzlG/EK1TZxVF+xhEH/mv5JuDMSThYf0Km/
M93MyKPYiekvI9B8GP3rcrnFSOCzVY/anYDiN+5NhEFhbKGNRh1wozlOi8cBCoJBUZk4jpq/0nYE
QgAKlaUFDkTlORSw4kF3zLfLNAurhwN3PttWm92Gze+hkRoAOlZ75VMHjugIo9OSj2RPCJ3cQLAx
4qelzo6ItsD1rSSaTDSBccsN0RNX/bSbTh3q1mN2P4WGZNUX/tscFyVmy/yo+bSTjW4w9q5fK4Gx
UJPXmVN8nKTjUR8OKYimcPg+RtovigYU1Fn8ts9EL9pWd05eZPHGddPfoQ7kPo3VQvBJTXXkmpRe
hP6PQUWpCG01YYvGNo9dboPO7HCUBJugApcaxhmhUPp5eT7BippQqo8uTCRmz8nHIREs9emg5Y6T
fp4J2LY0yi74Hu0EGVdYXmVaXYqE1m3Bqt5LERfkf7w3T++y1cBZVj1pA1G17fK8yEbCn6WEzQhN
5vDBQzdqbdNf+4h1P8WhUeGzuN13E8xTdKVZ3U5t1OaOJmbqBtuEv6Gx3tcsxGXT19IpCnNIoWeL
jHzG5rDajsBdysyfGXljETqxCpUCK5q9ps5sBoFFBCTTiJ/Kz0xN0NBQd7glo11pQliIRzm9bdFZ
oLJHZiCRGpfv0EI+Lpy/7IXzSP5s9Dk7rdM4qRdCxRlyphccta8jSxFChCyBKtdTRx48QYt2Cnsm
8BBtGv/HqrR9zz3Pm/yq7Tl7ENmZ85sGMPjhp7rxaZqQ+C8am/x4PD1KxxpPQhRpHAGCrA0MRsPp
CtUSdVrlYvj5Gm6JIJsQ3t5TXwZdDT2hk3edl3mwd1tXfiR7QNBytdjH5WVA9MqWqKjYpEB9kaGt
QRdgy3qopttDDv2b1bQbBGR7mJi0UCr2hTyPbOcK1LGEb1y38OYVIqAePluEAbMjPBMioZsJnKDP
KRlX5Mvccjl2oV8tyI+AbWYfjfxUIKqtmVHWDhtzEPTTFKAsGFtp7zToiIaMDLfLGdXf711Dznxc
GIv5yZADbvg00Bt/1KbnoItAlAhpYm/s2N1wOOg+zpF3Z3KbmaaHzmrOn/aXMgM/O6v8ItmfV/0/
ron7E7QJJ4v5ynFjdP8MYS9cY2237VyKNVG7W3rHJUPCkL2TUWkL7RUZllZX1Tk4gK7hINwO88JM
WBqf1jA8GDMtADtxiJjyUZWqE7jlQ4EomYgHscIUbUPbwoyUm4h29oCWxJcEwiXA8LCCEeReHa27
REr8JVq0KAFm+pa7TBRIweilzY/r+fpkeznEAS4/wLA4b3t154lalO2sXZreLas9M8ft+uZmDi1A
+XTPP/O9CQKPVVkS0ze9RUMRCbxeMBf2SavJRshBL8on0K+pVmIm5TE+c/JVZRwbkeS3ItP+EH4f
P+I/o3bIPHktEde4EYuc8r6TLiNbso/qNufg3h9+BHzIkMTlk62ZZbseaYHdYDjqi9xjMvH8OCTQ
t9VZe53IHkYdO8BXbnFPrhGS4YRH+UN+/e95eGTmC0hJzFppbZ7qWqviGWlLJwGH+YUAoyXn9nMK
oQSQ62WX4H5M8K58mciSW2sA3THQnW+6qlbjajd0WETazT/LBZ04SVkdA/JPN8yfXYilB/9nmByQ
/H4QK/96301BaZ/de2SEvyii9v+6YncvIrnHDwKY3l60siEoiQ5K+HRmddaG6wiygwhe86FGEC8s
mcdXqtQQlFYSCJcsIemoGDFua/w02vXez+gfewFDV16Mws16R6V/2U9pD8m1zx2VXrpe2D6smFbl
6g+CSZM8rqgoh/BlaSj2PQ+p9PkRwSORsZgXeRzk7Vtd3silVU/82HcRR2XrQQuQ0msqW7CIaur7
9f5l5OvRCdiCn1LBVlyAWy2ziJU2pclHFrb4oCpg+7QDsRubJZncIxUfM8cRbbZd0DNsh6JlMku1
wQStHVeJo/IwQfaTu63LjDsxCYsvAN3M2lLZ5mhzciFhzE56CeRHqsAbE3E0lIjHlieXucpxXuSp
/DSIL8Ju9JppvENCUDE6T3k+kvSh04vQ+Igd5oYcarfXddkKsjMIHEwo6T2xHI9Vbg6TjUmCUHKH
B8DAJWaiqydNaOEfVe4RR1lvNKmspxxJTbakbXUypfJD3AWfRFVkRFl0R8/vOaUt1lf56JaBwuab
jmJWMuqvt5vu6lhqHsal6IrDTXpq1GywK0rGoWpxqy+uLNPZ0B053fWmWrDHqlrFTi1QOTdnrmDR
6PIKzsmAYnD9eja4sQ9eujrnp49JeBGdNg2J/VT1SF8Za7molYb1wrbi5QONXNjT8UJOPGTsFtKS
2ujSIQtnCuNtwOZepMe+kLF87fMjvFT1tzBWye/V9kvywkiHOX54BgBvtvBJnbwvFDhRQ5wQyw0F
ad9SXPde8nFNJHf2EZYiYAQWx4FroZr1v3voWtYDKEbzXq/80jQTUfa7S7FDi9dQ7A+LBaRfTsXB
VhI+aMWN+y+D3XqZRZU0/c+YE8HbO3g+nCagxD8X9lR5qDVprvSh4muh53ls5ZucLDZ0SbmTEfWA
LKoZJYNVAKOQEC80EoHP7K8A+h0ufZ0FhMyPhHTDxlmITTdeGj8g8pXw0WAsYoMvqPkydRR3oDYQ
DKF43l8/ULRXSzigFtEMhqXxXFlbF91Cb2V4LcmGtUB7RYiB8i95ZXvNam0AXP1H8WjB+jIJuYnG
qJVoZbSYl7vGyKuW97QplKxzGaxGg7hd/IoODpRAa52hrWYAec809pfGYF6lRTr7xsd1BQ7VzPbV
jI/YdlddeH6PdFSY+NqWr2Zq7VqNHA61cR24cPc6t+qNoXZxTsT1Yym7d+6ZQGKqQtY4g/BTfm45
rZHwAsYgOt5s3xx3bf1I3TEPJKsA61GvOErjWCNlIJ4YnR4KToHtYVV+dhNAaNt8L4L4vKB5zxYb
JOzSu3hZJfYDSi8Aj8vJ+oPHA/83DdPpBAZ58odhPI8Zt7AAoRxc7Oua3DqbEpjp1yRgWFie8zTn
dT9KvRuGE5B/mGAyFLnaFwzCHL6sNtPW0k/dsVhyMXx1qe3hhyrCBNwWmKJXGKgDHWpjYJ+kvsmN
TDjr5GdFTzz9wn47uX0+gOwT2zNp8OzT+i9by1XlIpktvfTbyQNQk8vKT6/XBrJ4UmBdFzucgBgb
ct3oONJkrVKhdJCDedlrgZrfk3PFU+2Dc0ztN2TsUJoKIohxJ7k1HEqHXmyhIXgIyJ6ECwqYHPTI
LeJf7EGPCHXoSVxM9tuQzXMchsOCbD+p4JD5AKQkKFVfYFVrBO1BdaAh7TH0vqjI1RwTSfF+Eqob
CxIb4/fQ7to8FPJ0OBFbqceU81E5NJsy8q687qOVP02w8jDfDztd5NH7uYDBYgEtPIGqq6SV6loA
f6MrGRA6nJO4J0DLlb4vNBuMa2Y158G2/TkYMjYrI5+pv0d/GXFNvO7kfGyZAomfyO1DIa4LePbj
OQA4iapEm1D7+r4cZnea/Ed88fL2wxOZj4/gywdGb2GClHGQBlocsvNSlVijtPiklXzWCM6TMvly
E3lQjJuss1RZruBUiTm/5vC5MQug74Xl+gQnqJODmcqH0uQqMm1shOEYsqBHIx2WP2r5e7S0fkVI
lZiGsRO7hUdmDIEJaN8e4NHMaYHYh6KGAYC0FLz/tWzyqpGfQtaJ/nErQSmtzUPeA18/SrpXGj5J
TAPN2v7gyiZwAuy6QeJdFIEi9KsqjwZB2lY7XwJWe5qp3+seQ5UuPRDfNiQ7Lw+M5Me7Nd8P+b2I
S/MMOJtXyS02v1kVN+I1/epeY06JLE5j5tYiLtPZrfQx8le1a8Bvu+Ymr80qUpme9WVLZCBbQFHv
S/5SjpjMOukoi6aqLVBb2TdlDx6267bV+N9mZ26+9RLCcPOg6D/7k6A8vRuCekUcdNLZswumaqkX
WngNmth4jRMZXhqSThFiaQ6dA0CODaO0OBCB78fK0mwezpxigQh3UfBXhXDEHgUih/QAjaBSGhik
Zr8pCmeLwSgd/MAOHujhV9tSS1Jnoh+EdD27I61P71lFFY+n8NA5tRFyY3fbI+HDLYIRbzHPAQ1N
CwCGSB5GTUIJbczfa1C8CVc3TfwiwoLhvDpoTWCld5J34gG7v3C/L/wWw1UQV/1OjrDaWUGiodWs
cYX1Sv0GPn619YC5pwkhOSvzrHe08GiKUQmqUoeucIjn2VgUKd4A4G+MT4X4vfnF6RyAbf0LsBK6
PecNgV4LUXe8QqReyjP3u/awF+uBFHNnz/FPkHJHdREV2tUSQfX2sdcCTuoBbFTmHxlkCKi9LLZ/
YaQezxaMMIDusPWM/Xzt52reINYfaOMMn0yewglMMcaH+jUP6S3lcaZXu4VSIn2fzZibYPb69CIP
7E+KLJilGqbAYgkTe59wKFfu9BcT4O8rsve0O8CYwrG5Af9I9UijtRarLfN5j5sNCX2t5ejTXVj9
e9qjq7hHuAaP0VkrSbKeSFUosWcxYwqlee+PQdANRmWMDE9aVNGmri4KqTZw5Ukeh5zbMBMy2Dze
xIRiqh2+sbuSCmZklCDe4vcHtGePGns5xHE8H2EGSQ54nW1OoFBxStWfPJpLJDsqlQukBxOEEcpb
DUCgcXRJGLlfzj/YIiracUIL6ECaKt5mf+gxpIybjhAq8gg+E0/NNoqIy8fmckUymSS2BcwS1LlQ
ZzdHXZCXSWXQgHQ3MD9yZhcbsAhk8ys9/2Z1rx64WsdNxzAtqTi5cMyOf0AuGpF+Nwej597r99X0
3J8hrzWk8SasqnI1p0Iv4bLFOgetzoH1UDxrO4YutGSFK5QJ8DFi7X8IBVwUDCsPw2/4LYjFjqV4
QocpiBBxH6j2z4qrqdGnxYzDuMWu/hGIVMX2bY38DCfOVZXphYR0HfNM55ezG5XtaLGO9+VBI73o
ROnAOBrMefRjC+INZ632TDwZ6SXbrJXBKO9uTZ3IqcDivIotBxS/LkSPI6yqm7DD+Y0T2Xz5QYDk
84L7y1TIbfP3KJIEWRxkBbiObwszsescAkKMdnF1EIKDJ8PPREsh2NQ5SjS+HD5i+nA8UmZ2JS5Z
iTYlLOZNeRMqp3Mu0l6LdL5L4sranz7QmVmGOgTgWORjD6vlVY5AMB8Gc8GdUSZRTFs3CKYd2Bc7
IjRWYm2CPs+7jdv22nAvv8NAeMHxbsWP8qFzGvkPV4ySiKcqXZMMZXvKvkOm+g2l303axoHYzvl2
Q4IZztTMsdWwn/WvPxwNU4jgbna4pf1QKwkVf34YO9ux2p9n6CgACD3ZuJadLwMP2DQKS4fS4lMa
2uOZxCY94agxLLn5F0C+Uxd8uHKMMzTLgeDylUAbKROSzhLl5L/rJtkbt/sMlSjbWV6kexKtcERQ
nnVkKn7FrCL8puQSfjQc6uNUBSI6S072kzQvapU2fWULZo5U0dW14zZ2ySavhBzJMAlZfjHgC8Hd
9IamG3cmT4GK/GaSSvOaptsMl9Z7sQclubisXVZ1R24oPDuwhYwr05jfGJv/qF+JMvB+7hpBaWSh
rRDgF+WXKL7fyIyzDPRiYcXcWJTKdpS20t8B9H37yVBp8k33LA1uDUIjYA6t/+O1W/66ml6H0uza
sdC595zDc7l+eLNey3a4p4YDousT5iZ/UuI8S1D/VGpVR5RJSX5YIJzuppBv8p10W+z9WbXMuqgS
zGFbhXRIVyFWlaFzuobJz7yWgtNs3jWwZKe8X5CQUU/2IoOp11lPwN1L0KPuM045liDNvXuK+jJ1
L2TeKtO5vv5u0PDEDQnLyGh2sssDtvUhQK7D5j2kIx8KriZs0FLOIifTpiZhvPoHeG7NdKN0AL1D
0yeY+JW+JaG5uw6S93ulTZW3EPIUJ2t7y4OX0lLeLtNYf9vqqzJg3gkWh2/Lt+AdKo1qBU7wmnqU
5Acl8khDbkZP4XSb63RzPFiQ4aqzSjyrzsQlFNjLnelyaG5ngZgiAuMWOtTgjkouhszAKHVJ4PVR
e6BPCcSf1g9z1k6+Zv9UIX023LFINMwQvmGYdME9h5uLoYi38pRA09caCBEbg/KcC1eItVN8gBKl
lM8BZilaZxe2yozhzbpzNWvu1/w+Kg9hQrWXnMkjhPYg2Oy5A+lHIVYra/OcJ4Se2hH8oRC1EyTp
6rr3ytDfUlL9Bc4WyGFFDiThu07GiNnyjIpfeeX9FV4LZfcnbEz5/5tgtO3GQZLZCb8gKE6gW79m
aOWhhzQ+iV2emaVrqAQqI4ItF2B5zIlmAwlpyDsF3rdxMbe6oI5qE/+FUdLb7Cl8oEuoJSyXRP0i
5GXPdcax5gkYF7TCoEhKwoyT6e0Yaqrg3IyDsXl57KzhT5g6ihAlg4W6Kb+L6ozbnRbjWNS9r5f9
oUxh29Gj3srcE1MLGE1+dlm3aAxhMQMY1eQIMc+ud0hyI4iY/PeN8UXRpjmCXhXxwRYimmGVro+1
rmCwkvOZtNC1Mn0g3zLIdSO+fxz2iEYM2mdjlS1i58cu9p434F78YAWeyeU7J+lRnUMNIBa6Zj5X
ZH012rfZJG8bRUQUS0oniUjiZaJ8EWlBcb0dZvjTD1VW023BtogXIphrbtRbSFohfvoa3oGITRYi
ELM6qND3vkDAHRTsqpJlhz3mOs7PqrEnj5e0vFfFmb+K53ZGzoiMQKVPoehmgrhoOCwSszFzZocb
w1sapBz/2CQCDv28eAxrcQPObMaMdPFghW13kgE4ZmNybNrun0CBjwWXcoI0JWmmjfibtZOWBcx1
RRAdO4/Mt8RAwsKJiZ1PoJYfnk5YcgyC9qUqWpUBFIa7ceqyTCKwAfNnJatSmbfXb1rpsFK4sJfD
h+1fXUU5bAkdK/1HORfaQtcsKyW98RrGpEjm8ujFY0UA8hzOAwYpzez5vXPVGSC1BbD1aQCo5wkf
wZpY+T+KB0jsvA8vqMD0AGWSdH5yxAsTA0NsK3ERyGeZ9HCZQLqRHdDioTFfmoLAc0elvptwAp57
9NIdVhFWy+6IdnTmIs9/sHin+bmzQN4PAeDcIemUocLmGJotA8tb5YW1zNYkx5x4epr9D/vCIeVf
T+XFs0Fflcz8c2IPudJIUOXkqFH+IIszkIU900TYRiqlC4/mZ8WswXw42f7c2+p6Aus7XJceZAat
0mVBguZopidxvltFlRtTUGNHd14xHvtW22yZeKFVWibpWuWUjkMaDT1Z80RQ8qDMLSuPGezKxaAW
JYHM7VaKcUyt4takOfQYhXpGMO6GQfmS0iZYVkPgj80u6KmaHiMPFtDhJmt/Z/Cly7QQRqJh5+Gv
tzbu6cyHIa3uNlL4sF+KYcLIIX3R/0apVRJU7PIrRqwc9G7sb2Bj1u355saNV2Q0jcZCdyshyugx
UQJ/GhT6DXzANuesggbbc30fMEFZ8lvk5ar2w1rC0xiLKTbtj8Gja4tc2c5xP/SJ5XjQyTvaVoJ1
Iv08n2v4f65TNNQBmtcrHI8hw11hChRsDxWiN0xHNVaUhNb3oVB7o2KSOFbkYf4jiY35KvTQpskS
3n/i0yZgcS3lUY+bvCB0F4Kv6K/Lphy5RTP9K98OXqMQq661omVOq4QkErS1oQ5iive9fActz7xD
Zakox0dVdcCQ3lLhzO1luy3jHIxPcFYRjBiuscohO5iV1vwxWEr7BqFoyQCzvAa50jSxfCEDtGAw
XLJmFjSEq63iizE1QJ5tYBDHf5bpplkSb4s9dNO4z/zlJcE695YgVnlUVIjG2MVilh1KFPtmKC8s
VhEQ/5No5VZZGkFjaQwxLl/N38P57xSQW6SfZbRMB0ta9PxtIaJocseaVCMvhelR52EhuS12MjZb
OVkIzH3uPcTWMLl+hNBMp0ZLsLPloqrO0ZEtqF5HkGSGMOZH/KAB/Sss2O1uZpgqsbLvr/B78uIQ
IJul/sdrqo8i/9iBh43+Vurevl02Rc5VpYfDsIlXVLOOHOLw0gfflX+rLB/h/qAxBss3tGu4xdCT
5trZZAetft+LijKY9GdzvU9h5/2C6UAiBtX8A7l9J/C3nWVsB+zbHNJ5HS1hEsezrSSWLZnvIqvU
pJyttLaJrgAPJAHzKo5fRNPSiZUtNGwHhWwdEE+FF1Ge+kjn4/YfXRWOg1wpjt6zY9Sv8cN2gwKm
pImJWx+1MngqEvfTc3E4cTFlMVQ/0/h9wtwjOQgm/tR8lFFCre9r8vxCX36p6dB8R6Nzl/ZGi/I1
ZGBsVzhLC+NDKBdQJDHSMCaBMbidulrN3Ng/2wlyup38dKCsWK2PMVx+Jrc+0hGF23AyiqlislNk
9MHME6uthkwVrYpEaE+sWqMGWl43wvnAjNJ/V26SIWKzAWrHI7QZ5JqhKKWQgJRK9xqU4kaLwIwc
3LVGih4QWArsTfN7xBFNTDpWBtVxaaRR3zfrh6LESfSysC0itLdmRiUyiGmdUBnHz3M7TiBz6qZ/
YOgUWx36DuMeiGlTfFMguhZtouf/nocT1sy1JJIonAjEmda235A6MXxaxyVIO0YTeBgD4+Y8fWwP
/HFaNhwp5Ic0C6froWY4U1Xn9lKnstrcNLAD3E6F+tAs3n1vz5uXuVgyGcjn9oSSQvi7V0ZBeK8w
8R9sESpak1KM620sWLw9+rtrTNHmFGL2tMm7OrLxLqOkUt4GYTLUZWHdNZIdflTAy6kiRHh9F9sF
PyQlhaGo32SuO2yZzYMoY9YdRdymfrh0P11YZE1YjRmBam7KgfWhHUULBEI+1cebH07Cu232stcj
NsiVcsaR+b6nQ4o0B//yk2w9Brh4XilfQGH0lfFzTXhQUwxY+5KT0F7xPTUQa9ZEtwoUPYJtDQbb
IRaHoeO4o5JWfe5mRsYmvy7VwFV7zXaGLILopQb12aNPV51SbCPoSNBFjZzYJnGGdmOimheh7RY3
cwIaSoA4V9W/bYhN3OBWN+nrpcUie3nmxQplzdUMQAmwh6xxV07lN3GtyraiPWj1jOnqs35uHXfQ
TcqrN4HHOY/HWVwUUBm4jguZWPxQVBqscf4+4e/zjLE7Nd4/+JoiV10xA/16selLzGW5TeRw2Dma
UeLo7aSYCtTSOAwfrYzctzfnnSyjHVML+L5uwbm3jOgSMAAxESrT1cWOSrVgSOTTLh7wSMpxW3uq
RZhxY0RQ9oHmTrXVYkXIbQLDj+KXeovDFnX93Qz1BDA3JDz1ttAqFXauusTO3or85ZDLyBbLD/in
Qs4+07y2dcT8PVYKf5E/bAzR72bj5GK6ROvXSoNmIZVBys7vml7A7uGU4d0dC0o9o9ktAllt4yY7
aAG3U0CS+jK1/Co/3UKfpsZ7FMvCqz8oMDyxo1V8LzKF8OatGXJI08RtyUYKSqTiXq994hrOYdDJ
VVGsHuiyS7tPtXixwi1JS+YbHNiBvp67pLmqCCrqVIFl5HhJFa+PTu4H51/b7OZun8/dXxcU0aCq
+QUQSnSsV3fTP30PNe2h9Q4ekSP/v2Pws2cSjMm4Y0ecFYqAzavtc1bZhXqW+Uj99WybcwzDd9dh
Jhgl9hBas5P4kdicLL1FDNe1Uvo15wdFDnw0owvvoWtRINVWfdHpps5zcCVT99xVkOHBTf+L9cst
oyJPJMfgLkpFmTCNocKX0xCRGhKkZAGDydJOyiZOnmbrAA1PRORr4kr50gFbj1CN8WplY1VTko1n
kAUBIiuDEHNWbFsuJ1BDhca5YBaSrdkkz8DJVCwLOJ0z6s5uA9QUcJUn9+OB0GI2/pP9nhJIJThQ
CVg67vKeK65cJou8dDO1ORLHYMMT5xLG3vJq6llz9i0Z7ihdmjcKu2NPit1ynHA73aCI5aEDiRp3
jrabAzm4tlb0Uv5nzpZ+xpG8YbRKypPjUqgaHqX4neYjobPlG9RbjbVZh3KGqOi/DcRgoEgxpMFh
XjKXpXagfbF6qXMeh8iXaAktmn3Hd0QnDijOpxupQc+8PGSMGqB7A1S5p1Pxouc7/b2t27BJLQPm
RpAJohFGvjBsM+jvcsR9nnIpTJIML4gJaWMxbiD1tRxHFmMqhSYYFbhibWtdkMUzV8bSyi511OBr
jB3qzeoJKaO20Ju6yqk2dLd05hDLjrHNsMQfp451ETIwo1ISylIWnf4aM96gsrf3v6LJMx+pLGR6
Jze3cMxlav9BKM8G/ZW0Rqb94HVI+nCox+GUPx/Wj+LHU9z+i8/JjRt3lM+S9ETFfenDWXo8TA6/
owm0hOmOIUJDfBOGOjp7X1OQcz7VXnVV2jUr33MM961LrfJ9Maj0ph0EIhdyxf3+ah0JCGSCz5B6
m2bN5D19esnhAivUyIPulv/3rKzhX2QWHKeIeFFU40gsAHv+P2qcW0MkPDa1ZY480iMhT1gdvl+t
Hp/lKNHBpTozoYR9Od5HKs57bfQ4bZVBmGLDiGmsfxU6v5FUXutFWyDxSRja0ik8yGWhmuu19Apw
RpPWL4bNun9K0f8vc3xuR+RUEWgkMqFB7OcJZNTzk2/hevFEG4ce0dsbU0gOfwyYlAM/AwII5CWM
+3poCpPR1Nv+yWagSdshzqzaTQ+dbVmUeUyc699CZvQSi0p2JnGiPKhWQbqYZ0S4hzJWAhyEbze3
r1YFAU0g+4oAR5/kosrDeA2cHa7cL/uiuoe8TcJg46wYVf73sQvR4+51dEN5fdhWW3fJQ69i39Vf
NdogdEGEcgLpcDlLzO0axwO4XoqFUCq1jBuiMjuFpq/wAw7U4khBIYZLmMB+VNlG8oz19ekT//U9
fOSumqaKuHrehB/luS6BALC/VZ1tGyj1yRwi8V6sim8YzGBne/GpJhgL2l1l3aMX+U9cPTli3qCD
p8LVkIbtBD1+i0UD9rwg7crMNulgD5fl3U9NmdlVGJUpyxIITJDZE+3z+tGaZkpLqaUXLjs09VFA
fvRtRHmktd0g4cqmPQvm0Emxxe7lyrSnF7i3b2IGAoDbI25gP9nHzAjlm+iruT4jXbIun3RPwVEp
P95cfjugLgW/GpRzxhHGEbNNarmZA/neEnZ98iPb96LYqT4bodQubHK9ktdLzGZAd/zRui6F3L31
Cj6qa5ZA4hWZZrxYjveHxXpqi/0RgJ59FDBfdNbkmlLdU9tLbh+s2WzxROO6W9FxkCPkDEBDnYhL
iIuQxFgFwnkQ7YVl+osLWOTXdtdOA/K/jmJGtqBOLaAQ2/dmYK8rwX3Bmn0EQmNa//OJDZO3qNBq
0UzCNWilMVmLJS4WsqWXhAp/cv70ccJfZLsQginT7aO6YBi3JhTTqbr71aUJvObCyWLW6tsmF3iX
k8URhWfFgg1r2XjhnCf6X8VymLQjHnTkkIBQpAL54DmqeFocF63RxR0cVUmbIg2ZuPJMOOCniFVz
lPEeCANh+/Gx/atoxvM8c6IDE2cwMtolKaAbBwtj/LMBPTmAdltyNGa3FICMl0rFKIsr/Z2roN8a
yq0H4zgeOlKJlL13wQQAv1lw5hPEcHX46SnKUZLOFlQy51xl/826jFgG0Q3Ig1P+68h1Mqs55Krw
tvCmpNPZOxGsxwg9XtSD3UcLBtU5spHe8Cv0XcmyXmxN00stUQtWT4UCJyJUUsnChB9ThTBR/FAL
0v5WUI94JMBhxwFd96CVJ/uWaS/46VFDfMfdznDdPkOGZouQQvpFm4LnEZlgH3onxw2pjdRB6jsN
SdLktyCRb4Cb1OTKRUo3otA9UdCvkSoZjRCqBmKHDqlxu9a8r6wcWrgD0qvGTuDL7UYTxpk0bn/q
YW04GMw1Ua09nhLzXojz4XfnQoR34JS2HpS6/T9Z93956iFGqPFlkJ8d/3N5MQMduYhOLxwO3o0o
OA72ahc59Us4pEKnJGI1NOtCZh6kKFRjZxNWHI81mx8L6RAvCGJB5LwxZJjia/ASEJMZutbqz7vr
ojp0dEN4ibT6B/E5aU33d3IKB8vBzYQstMTRUpq/BfXRNxnciIu9Kjj+vWmXoytKbnpNOQNDd0Yy
ewg0Ip6z15StSVEOvMgnDy7pZef1ac4KBfUZ2qJE8Hq+kiduDQPQUIN/p5dOCV7HzMLXaBPbRj3n
+jfZZxOzpr2or+3S9MIOY49o4q/l4TeIGvtRFJL8TVCxPWrxbmHZaCU9L8A04YP8c2xDavab+2GV
cGW6tTaCLGyJTYtB5jZecaxX+jBocUI3lyMApqK6kUWUNZ3PB1j2Pf20a1AqcB56lD87+kW2q4YT
GyZj63JQmHPkyOrrOHK6jAndJiNSPvPqF5aBgX/eo5WJAh8+z2w5ofA6DI4ubi66fTas+i0NRXbm
9uIJcX7J9jO905MJpej2rXLNsSHboGd+EB9Bt9N5OOX5TtbyLjAPGVaMfZvSTn8b8SWEVtEFZsYu
LIMwrbPX7+HasNygJhNicLBfuPmtErl+8JOUkbG7tPLCZBt3b2C422Xeh48dyJX4LhsAJ4XzhKig
GMAvm2ey+FTgTh6rtLOjIF+TEhx7uUB0fVqIUJ6XqqorcrYvkGoRm8GdgPxTOq0D/KDhLOlT29qc
/2Bjbz3NFwoUYPGswFhpNU+bv2tVh20HT8Z71lPT3h+RADqUySALbs8nWOqM5As4jd4Zd56DSQ7J
5TrDehgjn34Fbm77adTDM+AnwsGoBwxyW2WZ4ptG0jy8l8MPfWQ7L+Uk0gFtg//KrBYvPgH0Dqfr
AKHOiGFag5NHicbYia38p/GHsHI6mCaiwIx0mwYhJTQgEHAxQCL0nj2tlS7i2tCDdhMzlqcdoVOv
QbsuuuQJj56V6hK3Li1mLT9GE4LXjsXYRDFv7QSu2jkUuvZ8ocU55OUiGmhf8c16R5cYLeKdXHar
/WEQdRQ8aoYSm4yTcLCIKCHWdU+PkafNrV1k2vqazQjW43Si5anmxp3q3YRpUb3RdvJ2yTdp72W+
E/C2jeplkvOpZRHgf3OKeYYsH+S+erC4v1+Dd5DFBnm+Q3PSq8N+D5CLOnJ94oxgN7nuB+QJuAji
ZIZXXHCCmqskPmGYOvXxvq9420/0DDs8cUxL2iO+5GX+pXfSoPguU9ZMSoPrPxPeuCQFZl6qFIJH
k3tZ7qBaBJzFh5FES7AEhC4JNPsgAaBzc98y4e0ZVprStFTfHD0dumGRqHt/px9QvvIkxrNkL/rD
fXK5BC5rZC1qofx+T+qO2HS8WBVe5KTcy0P7g/EuSfu3tcfUs1+cCQgRilSuTL+5EBZC1zt8By0+
JmmsHrKk+L5KmGlQTA5evQVZ7YBRgGAJzeFXAvcuRn26V0zUHuXHNCuuTxxLOeLsCsDyFKG4lfqZ
HONttD6O/WCLBjM4Vff3mjYYqAlRuYzvssbg6z/MVnkdQfRAqIz7n1p5P9vOEU3HaixnSV2ib1sM
vrLBt5iUZqBRApEH2DBBHqzQ6JrV2F/w9h2U2/Gv1BAtzVryzxnuhmlUkMxYbNmpb/W1PRHit+YK
Vd88LTMBw1LOASLOfKPi3EzexwjDkqdTkcqVP7XORGKsMdlCHxzAxGYpEUbvYKCZ7bZjwqJ+wWMs
yr59egeQtceSy1ITUnEPlJ7DrNIa7dA3de/8iWq5xSGpOF9h3phj8H38c7WLPSMjtJjRmcLk04VI
ZD7PUfgKsMpQSiLmNtNNwUm7YjYgyRLoejqFeb9vgagMFEjq+StFW93312w2JXmnwstj/mrOhXv9
vjr11R/ZeqWzL+ups19LNQlGukiQl+VtOp7yHJxz2xuAUQBcjUJO4TI5WQqyKgybsZcU8khgaktU
BYqSyJ+734iiSqAdE3K5aTR/bnOL45BrQDcjyCNXz5oVAF/fnbp7WKASA29eiCeTeLYrX50qatCH
I7tIgMPHPqmGyD4ElOebJVHE8bPZRNDcJP/EOCItsSSCUxYiBygXiFTmW06INmGiG7Q9v8Drf77y
E9fA/PpjRpSxhjj2BcptnUx7LfPn7XN/xEXA+cd+uxBSmGx9ccARjCpXQ93yRRgbXz8iAHbY9Ip+
p5NQI2/iukY5Id9QfeLUJ8YIg3yKiJNCnEH3hMBlcczE/K0dy4RpDrHwhV1sk6mnfRzqxwr2I5UR
5K3MToQ6RojjcHc9P0Du1UvuDfJTdYNHmru8/n0NrU/XswmfVdg7R+LsmjBNy+F+29/IcGdBcrIC
bubWd6FwZYJ371vJfpSyVBlvY31XTbMpld8SO+6PAdu6i8nObMkH6T/zAffM2xEo0JIG34EwSmnB
K7gTt1qRLF4QYVn9EsI4AxChRB6aaFqUK7tXkZDvvPexmckEZqcBGfN9mNXTcVNYlOgl8fUvu9GV
kzsZ379j8eh4HOz0ep49suqGz6gRC1S4JrcXF6ulxLxtcc7FAv3OvSqd8vmSSGQCvySIlEV0R7dh
eXYqw2y+BItU0Wx7WaVkpgHrZbShhbykPUhWf1gougra03D2yS24HquwE6QWVtVhZ74FxFdTthyf
fH7/T0mcWDpBiZ+lxSsFZpXdu7yHUuxrmFoE5F4qCRcxyX1Z5BL8pVj4IWVJML/qKjbLcnEV2iDr
7N7sRKb/AmxUL/08va/bKbynYS8orn2oW7V+nIUAPqajeiFX/QZNJWxfFVpeCFESwSBygbeYO1vj
rlMewTI2GWpnaZ3su3Nef28QUU9oeqqHDVjkUb2QmNpopY99FE/NRe+ssprxp2iW/Bz+wFo5u7zu
cmQdNdtT8DgR0rDQWaa9VqBxvGu6GPOcJX5CWi4XeVsOojPIQxagQZ0cdJNMuCk4oPh3XeRBR7ZD
3qcsqFYNKR250SMb2hecRROu3+DapAjVkrqCHBN41nxFKNMZloqVGAMAnM/3ECxT5RaVFNnZF+Y6
782NgJkWKJzjxlqtva3Zz6hVWn+d6doUbDVORcremlETVNI4pU8RyHVcHNd+WbhCNP3M7gNyZ65w
IPKkAYWElUsXS74BPN4YJRyz0buQuWOjgUQm7u97FPalKcGIcxW9gXJyoFE/1CS0qlTBUVskECRv
5CgLjobDt70+5GZExHS/jb5ENNH82P4vZj0tokznCJULXMrj1BzE47LZoz+Sfs8p3XnV1QzeRjoT
Z6BRTZzPC5blWUBPhkr9DpqzAaLyX90qn+4Dv8Bw5DX/0CloYsV9j369uQgGS49iywezB03uwkTK
hrvzqEiA0wh7is2AXX8UzW8OifhdT10fVK67hIfLG/G3HSQVCgYBRP2dZAoZBHgwi1FP/v29kBIg
g2FUpmY6Aa3hTsVm5i9ucM+YCHBhjYvN+Zakzeknqmxo5N23HaMy3c+WrBjnhcmtEY2u/nLF/QMu
Ku5bDYiod3gx6Uj+oTspqbs//Jxs+1VIMZNqNF26Mrf3Xc1/REWgxJkjkSIlMo3b4UH1Qbpxzgj4
nn8stUvG81UdrMKTBbGgBMyj7DgfxZFYZf9j/vBj/egfrS0cKPwzZqBWiHp3wx2JRX0Z42g/GzUa
OShc97yjsPms48COeaS3EZ1IHlPZ3Ve/dUfJZZasqh3EvaMTdMhu5Mr7FMA/Rg5VnjCWLq3flwk2
JxhMc0lvlqyZjRiCkcCzZH7AuLAkgwvLCwfx3bqhFLHolpj3M+2VZbahiBI5nlp3nR1hTMsN38R5
dMb40boQmOfBLa8bIrdD9/HU24DpeNwWDY1r5/KZJut51fqTqUzarvNQ7z+nhfUqglHInAJbSwCD
SMrkFPDH98IW1fzhk/Dmxxv5JlOvQOZ2VP1u3csylKKP5aP/3zGsh8FCeIZQ6HkK4AEOQXJykB7g
v1c27RR56UJQ+JV1++G/47+S8YhBrL6SJ8pltDiLE3ZKG2tiIbH83HaO1lzoa68ddkYmo5ZPatH3
1Z5bUUejFeouiBTU+33rcV/MHbWDIO87eiEAKaG52xUMDsHwXVg5VCE6geVCUvXMWnvTtWULh2Ju
K6NoXWN2XGBLQTS9EGfkR3R3x9sgDtLmL5ytwEjnOSJ2OwOXsV9GuuzuObd/nM23tJa0+5B+eovu
LpEN/cuVFTyHLXyegzCwG0xRvTs2ONUZCt+k34Y3iXhnHJyTFe+GR60oX8P/76GsI5d6pnF26W41
fK5YRSOP2Jrnky4yCG7qHSwI0Gxuxc0B7Ndu4k0frvZtjrxDWvYsK/Wd+NcCJ/Bjj5wH5LeTmYwN
eBm7Q+JyPBB8RpFdhdjvmZRPbVdQbst4KRUJXqCxiixGMDEK3w79zTVeCKgpB42rDRZ6hSH6NePp
3gU1s9F3wgMADjg6aYubDz7evz/Gcf/yRCixXyFOkhjWLu8QdIWU8lBkjCuSvLqX5efN1tsPsLt1
ZaUknqgKSus/hKWCPMdMDRlJCcjaOEo9KM+qeaJSj6y7xplHb31rD+HmHMVImpkV4Z+BB1HDTj5K
WIh82eqdIaq4Tdt+Lwi6+y3mxyS5HmXq9ZiuPSmu28rSIwyp4TLkaAhNVzRvmyoKmvZyPaCCZ9EJ
duLTei6u7Yt/z59x5aJhsY+f3xyyYoTLqGncGW+MR7POpnB9gnV7i0Zw6GEfMCCpmZ+tzi2PzU+a
cHI3mTV88Q8UymOyvDcS9CZ2xXXJAOvl/rSJV6DUnM8Vwq+vLK8TIzKrFNoETSo9koTEnU87JPii
IuHGJc2EfKE3arCHW/j6pnTrMroOUDp4hLogJzwVVNGCmH3s+NH24SS59Q7pdJOIq0hKy+DOH49M
sevDFpD4IvWeL2xcixmJ1ooBRzd2T3IrTrGu7iz1GLFu/SH/B+Y6pQW6QjzSREvJUyLRFOhzCATU
D8r8GKlYWb6pLdwYHwfbSOVQeurt1mRCDIOXvNThYQqgsff2cIHcKuv91I2uyC77tIGDvhdBRXy1
4qEGtEoVsHdNzJaJnn4Oq9OxriUJHNRVBO5rOmuYoE0nmVk0TnPpVVs7C+tjUHaNpV+Gy57jcJkx
pO8ttAz6V23gjQvbGd+EW33tP57oFUWbFrdxqhbSiJyhbjSrLdeqMqRgTXh94kis41FGVRqdnLfu
Mx3aRQFfwYVioCrXoHUgZZzD9l2HIQvoeAUj13CbVjyxPHwljvZKh9ZfySqKPELY15g8Y4HUlZbC
dr7Let+vD0d1c1ZKgRJdBb5GSPpjF/AMjNlicseWlQSJXOcOSCmCP4ERpkWPENkF3kLHjF8PaIW3
QcsafRAA+dBx9gToRbsWqr1/GAgX0SFk6YKJwColBXroE1iKBPGnbUJE+VviL9BFQPYZaSfPZRYa
xR91ntMf2gpx4gozL/0S0xjOxHIo271vGrT/fxxhr6CHOvw4Z95vdf76+3QK8CwuZF9tyGbdPhDw
zSK/yQWjDCwT+Zwdzw3DZik7F+XwIaQUrrxVd2SUVyHZeKnqONvFbggTY6LO7jZGq6Is0QKXbgp2
nq9KDCtQC3AVRSmKHys6MfyusNomCwxdaaGrdN2Ky3IZvVhJhT4Vld6tpuso5heGxRkMouMTDtmm
wLXTNaV8XKSOWQeY81Ggk5o3vW9bnPCeosNh2Zb7zdmlvCLMfkC+fBGepHjJoIsgzAN+Bvlkapr+
Gqaej1lggUGo1DLHFLxcUIRGOEwnFL13LBR3ZVabyqDXSmJ0nntiaZnvUPbchQsHC0N1QTt8j7oU
6m2U9wmcDJjBu4i8lCXAHW/Cwea0nxBTDcGTByT4kx7Ws3rLB+lB/2TzzLsghqINYpj4QOf30PrL
FdWzJEK0CaBuSYSfAUAe9GRa60GRjY7Hub7gtVdKrBELECePx4IaT5CwjFAmCs32kabxbxzWJatw
UOEY3SH3nXXEQBJ06sN9cm+p7T1udZhUXdy+lScscqJs1z6bFLW57gJQ2GMPLWVIbOwjDXoeuQi7
s/wh+oMRR2nRpzcdQfS6YhHpCGiEXVISh+gSO/GMVdOyOQhaNC4As7sMLeMDiEJWlo8EB52cTB41
UatZM9l4KVB2yaC0YNRo04+oNyZG73mmIibrQWhzJZx3Z990Y1dVzBP3jeZVsjqq3nNCX5s18tpL
vvW229pmta8GmsEf4Mc6VbSDhyF+AjwLWJdPB0Mg9v1q9IgWkLCl35Wh2ItYo4nzhhv/i8sHZION
k1Gr8n60MasF2NB+sr8QkfsUogQVR8JEmn/0vxqql3SERkX0oYQkQSz0SS8rBsQ+QTYyufaiGMAQ
1wWwg+iRX6xjXCd3DDv/NqBWC0MH0zBYNx29+f3RDlizb7VwHttmMi317r3xc2YQUTd7epUEBxE8
+lXqGCYtBTIeT+tbzVE09Qn6k6UcknJrlE4hMP//q8p5KGRDpQKFt9cM/pZ39Snr2UzRWcDJSXbM
wdJNLtKN6vQRzMvvXLflBYnSPdRDCLK+BofQVghKr7a5xvgJioINaZxLq2S7E4Cia7/fRJ9NPEG5
+s5vkWzO0bipuQsmaJ46OnfVN9qIKxEeMHxZY71dtL60MDnx1wVixp/8zz4mtWYFVYt4B4zLABRW
bEvCdTyE33JLzpenoG/HPWIL/WYNwLcH773oFT6J9ZKTXXiErht/3UgeW5/FHjYQzvahx7zZz8mp
HWW7MWl38FpiG8ybTSL3021+2CbFPkklj7+Cjx02OeQA3DM3sYII/oSzRK6CZftoeRm3vnUgsKwY
eWfUnHjdvhxomgB+KSQnl4FHLrVzmkJJODHEWBs4776He13WhjHFIHzg1QslJUpJD7f2yntC3XFM
Wc9YIWlO4KfflRfrQg4RUenMPctcljewzso2zPgUFhNYK2tB1SI9R94Jj5p5mhHz1u6i6uXbvccI
iA3+wiVz7z6t7M3++M3B5uesqWjcSYRg1E8+Av8ImQ6dQMNHctLGYi1CWq830zyDAvLxtWDbsNVD
6e+hDt52g9FMGCHEGfsz763BBTaNLvTpE7LIDJk34gKRuxr44+SS1R0oaLFOppHslzuX2Xf3rUGV
3y2vDY9YxEifGMp7ybOfrcZQD6enboH2BhgcjQpvmLuo8Gz7/VZ1WI3SKgyVnbMFPgue7XHFD2qZ
Gmn8G2yRb07oBO+0a0nD7ynV0RBjl6HwUH2dDdoORA57Uyd8PKyWarBTGYWCubzZaq9SlU4XwxxP
agItizoRwe2AtkJ90K1P3Sn3CWtzoPDcwYS8JJx/e0dg/TJYPZmySnLPtvCmRCpyqYuDWtPh3j0J
1wx3cgSYSz6UVA4NpwCc3QG6lWyDoY2g25EsDcVhiOW4Sun2JtIBXqNej9mSwWiCBP3V1R8gMpJL
9Q+u9IXhIwl+Hoo5Y0U/sQ/LceHwz6RzeNpMmNPxGiItlFx09HgZuxHhlfeIypOlbaq72FWmQ75G
j6H6JoiBN2yVLsVb7fnahTLInQrVXMHm3hA7TsTRGssJDDfrM6hjabsl8jNTmz4k1LNAevj2jIMJ
ixcAcyrXqrgb1h7qhFXlgZwSZ/Kz23HZSInjBioKZ+kmQqtpDYI9Pgt+j54NPaq1gBGdzd3hLz4H
rGf1UipDwsU/WG7nIa9ubWducwJI8vZrUBhWaGO9laZf7f7XhggdWncCuZIGlHVxWV7Pp/+/b3RS
vi4lpBQt5ZoYMlpyOMqJ3TEkv96i+81qa76lPB1kmk8r0rw/QbOyiivwyz0CJ5zvBgSTCCe3t4/e
9kigWEsguloqui84RUgPsbfx30FiHQdZ2bboehPYE4lU0Y9OBQsuWeB90caJqI8mf4yza2HqnOhc
lrSy/RcZZsePkz4IbM1e34ny0IKoOzwtorGYbcnY+pv1HE11uP/nvU7g9ub85uNATac5D+OpEP+h
TzmOMiYWNq1h2a1vne3WYJtpOmg9oSHqbp7N/KJ/hxxPGEKfVWFzr4jEysfhgAPBd45FYUiGrWZx
4IdOaFzfooGcKqkuc2MGgOivioyFS6lEWW6EaTQ9Xgg9EktmacNMZlbwC8JnYGb7DbsMW1Ivl+HF
cXcGi+PPssXPZIJU67doZesGJ5ir4kpLpdKehrFBEHvNpOCpsyPl1WC9AWi0kjoZyxqE4U0WQGPU
sX0BD9mvhjaumuc47FEtNiUaUGBCT7LswJhdF6ACOZCaZ1xlBV7Gkh0hPfw7IpQ1s7tR1q5NO8m4
3S6wenhd1m5XbpAH0eFFO4hLZbMIPfp117XaYaTc/OblydxCuA5Qn8oTOJT32/cUqvwikEoSxaBV
hpquNzdjIivyC0g6PttCOV4hrUsPgjF0HFIMt0zOhLo6MT7Mm1LpDhMEitziVyyHZL13aq0Oijha
MCBMo8678iB9hPedDc4wXkFeHNxZJNUf3D8zhgjLzdDyJ74erMe/y+x8wAQrxH34jUCo4TUUJirH
5g4yPz18baJ84qk5yoTr/DRmSWvh/wlnVN2IukS6EVqT6OiGUrg19/rTzLwDBe2c0s/WPEmKcrbi
6lkBbgP6bQr+LERQed7oMz5V1PYSbdvyhO7vVF9oA22ysJmezf+tDcsukaavmpOrzoQkkjcuWxyi
eSRmGzBvYPIvkv67k086xwJY5/05ll8nZEfJg1nW5J4QwORDurEwJcxt9tZ2tebJlKG7dhDAWqFe
re007/yzKNMvhR714b5F1yuaPKS/n/F7EmRDPRn7v3cNugrW7BUaKAO3AWIDfZ2AgdFZXUChkHDN
djmCd7pAsL1n+1kbOPuWX+EIWsE7udAj0JNwSMomWYR3yowHwT0trRuSDliEzNF8d4DnqBNVZ7KW
Q82LFC2P3Kakv9pNYcWlUKliwT1yqoHR8l6tSwJiWCMemcsA0L0JlZHC8LNym++lDBRdgAW6gulH
KTiMSkXtmRk+pGBebCbjp3qFIUlNzx6LHCzBiPfF3sJGAVEzsIw21YPvMUxv3nnkmy6LqubC7OnC
I26vnF2L+QfAjfqSR258uBKOV4BeBoqYWnyxNKt2mFszX9/mycmIT+ddeqTZ28sNiMFraYMokHHM
crOlPT+6/IDU77r0AV+hIRTuzS/oqqC6IIWnl2JsXtfN8xQwoJsnS6oXHB7tlwTCic0KjzjO2Oqq
4STGnbYJhdULCF7wUkxqdfiUuMOor41V6AMRtCfZS1i6A2c3sIPLf99H8Q3ABJY31eg76XXs2386
oTLi9oTw3XyZpAhEPwiZqmRcHNQDyJdMbPYAD1h7mb2MAukFAmk3nZ0RmP4ywa7hXtTtJ4n+rTYf
mUldzgR298Ka6kvHiCrljcn+HgIOUr9iYEHNtRz3/ZGL0kZJIaZIJp7w6nm1qR1A3yMrbVcDo7qR
m8+lotXnvxLy9YUEj6SLQGpDCUWwtUUpHPiBNb0EU8TOsxDwxnbr48u1nXe/Nxbe52A7tWztyqaJ
sWrJilP78+WY3Jbgbh+SfCGME+O6CNqJaWX60pcFz4ynVtNAGH37U3KG6+se/+ucSZyhMVk/ik3l
K37EzYQuLJ2DpgkZtkbrpIDXG7yzr+uoUj4VCviXj2eMIwQZFTFppdtQw89kSCphITunSxig3uhv
dORI/KJKK80UKzI9ZSW+OYjxpRTVDWaWoLnoreVaoF7RI7UQZ4I6aIu6wwyGALlLn/MD6n1oK4Nf
K8oEAGDZuGAJk29yOpsb7ELYQSW9N0QIH4qYTSAOU3d1YQMz8EzY5fkfr1Ri2f/64OLaEDeMuHBz
JoSyQ5JXqm+dPQ7GtFh8PYUnqaly8aSdpyU27mTQjt9OAeb2Wxeom7QwLCuT/iEvethE9+LiveE/
byqyYIRG/Oxlmewnj0gweIQy3ZQDFh7vgePWEQwVNmO6ZQY4iSxx5hR7G9Nzr3YUMrvVXHnSKjP4
mJGjJiCvqZb/BbZN3eeAfjFXOISrAS/SPTmzZ60+fSjGTIwCf1z3RcMmhPR4RLzJ9IsXlj6Nd1+C
KgWWsL/mgxZgGWRjrk/w4YOFUPLYQm1vNdLBj1YzPclfG3O/zu9VeXNC9vq8ruGb9/oB4TxkJnfL
oTHPhSSL4W0Jd7pG5sXxZcaXvcYom2G6Hs9ELDbyFBWmxx4RyfnXw7CNIHC8JlKgAOZ3SZkZD6Zw
8CzZNF76c2YWXdt39uyMLg4suhOJjuDLml3/pIgILy+gj0hyi7HAKDXTI1f0/gFDWvoAmEWvulbK
TU5AWkuH3uVX/y/amHatbsHP8JXXazEQW72Ud0J4xcy+MbFpHXhz/DhzhD6kYEWFVR2fkIFTq00Y
OHij3dG34oz++dJWxKVuMnw4E4BKHbRRgrldB9do5SlM4A3yHjrM1NHgofkXBIrKtR4OS89Lla/a
wIEeqI/ADE7BRnr7R4bvshFJvakUdNJGys/CALETPA3Y4F+oMcDEG8EvvjzDsQImZQ16Hz+sYdHd
UHN+ycMpKsJQvB/HKgjjuU3j2y/yEAO0Op9yhOMPEGP/LkhmlvkYCYp5Tjyoy1N3oyTo/0E36hFB
peUGrvb9gyEkIRzX2tkcDXDZ/BijZYeUurtf2hgq+b7ZkUbmtRyPvd2Q3BbH/anR+bqfeWcpzeUS
bbadPKuXliyyfneSfM2mGrXPl9Qa5tI15tl6x+ueV3PWiY1palMfQQmmNgG9x45UKFQDJ1MVtTOi
nXCGl6N8AUQwuVD35xfA40KR11lFRnksz7Dlp+u7n/Tw2TQQmU91Y9Sni47MCLffb1Bh3xa1ICiV
qDVbFHaOB3GhqmCitPeJoZSEpW8Z/VrLHYgzdWjlY6IjYdXMT06LKc57xlIZWvwhzFVgpmokJuT3
eIZxSm+d9OiW1OFcWXV48MFDZ0wWCvaN2eedUA34CFbHrJ8fi0A75z1VykVkalI3D3rVd52RvH/9
s+EfffFYjFPuEpgjyOldRwiYOzIYbht/exCIFw0jeMfHKRPmeTvUMQvXRPCZXuaiEAdHpGRuFAc+
sTWt0211fCmkEh2b2/HvXQF9yAeImFvZWP1RW63PdYulUxmTokT/obnDEewUV0rxHJ8A1okstmBc
SuXKu7aw2/NoW2EkxFseeYd5AeIJwqqzfjNEb7g74IooX6pKVHvWmteNdoGvP1/dUTaLyv475ApZ
Gu7LirvI7Jmc6GHEoInNiwLePDO1vg5BSpmMoiIrxoIMNzLm4Yppn14JzWcPK7R6N5QKcfbD8amv
/3QOtAORFJydBHevGAewtuoZ1pmfGy5uRXVmWryAHOy8y2pKp5+H3ezX5BUK4o42Ip0u46pQS9oG
EQszRyX5kblGnGf9Gwm3J222eixRSRiKpNIFFBmHYANcVFdHzeDz9rQbHiGX7eylbvx+w5vuXhlC
WFRRiRu9FFq/fypdIVX826xO1UIdZBbH73G5zQ7z2EdNEb5hZ1ZJqoO5NOkb7ZJRpeBzUHUgwp9S
zDA5dXoiARZJT2AIONugWt8ZAlXwA0UScdO7CHH9SSp5A8l/3Q9dNU0K/2NWGUNk5pNblBzprADd
xceDqALVBOQe5v/2yzuIpXQOFhOiirq4Zc4EUB5vzwgZ4KMAXeilGerEwPLrkEPYJAsE7xxk1Y9F
2/OOhbAcp5hxjdR/E95VbemoIqEOXemQPWn0EAZwS309TVt6KsDNAMrluZ889dnvLN6oeLckh52R
ULFRa6imtPbB5v1Kb3RlASNCcvAmFJBFrbxBtobk/Gz5Znu/VbVe8Gr3CMpegyB95gJ+t4oaNbSv
KDmkrp37Dig04YOsu4wpH5uSFpXqbmexQUJQqTb/KMdST90jrWTMDhiocSK38nrzrQXJ1YCfxmhh
PRR/y3Q2xGXTmju3qLdqHJ22+8gNpa+2c6oflrPEFcLroShBGBlhujx91uJLYlq/ropprfXbFEz/
ZHBQ+0Vr6YEl0mIre6MU6wam/5rZS8Vis9UKqCc7bRQsIcWVdMM2XVY1Rmy0MZNZwyU/w72jj3mt
Gk17NxJig2Y92FeoQGCJMENcgwEnsZn+JQ81LxoY9tttd1oWKpEuIKM14CjGAnX6N4GSL8Bw5byB
4y+lPjaSdg8d2CD/Ud1/wq+6SmNC5Z0YSl06GUwNPSNk1k9WM8RFh2iGVLpwLofKGidMg8Bg3lZc
JHolF7UR/J6vw0fyI0p10BbXX6UoJzrR3X1vCUXarT2gR2gXOon6oYD+SLJGBhcmK0XsXotKlG8g
OsHAwO/0UnjsTUhhV5LQwnkWoRmwzTrZzRj15GXRkHsSjGNyGromFosopD3YTFl4uXwDMDxy+K+e
E+WiOkmCPhYczs0yU51wicLJEhUFglBoBWwaCgvKLZtmnT9U2+f5GMzzC7NEd3qhtXlUGgvOqEiV
kbm9syItnckp3JUif5nsvr4TFjlLkfIWoTjxq2RcziKnJ9Rzdr6Fz9hCesNMUQMmRnhTHxWZAvKS
A9n0JnY/qKJt+FbbcV3VdgEjTGT1ngzyVaop0eW7XneYWT3WCWiE65ebyIksepZ+/m4xpoAr+A0N
BIYrY+UQDzrikHDvbcJCnHkQQIJf8eusVZUgA7ov/jawlRopjWBRxqDmJePPpNCakicd9qi8eL4x
hRM6TJ1X7QNcH1iOmfeXH1telL4vGJxxe40ow01/6IK9sOW2DsiogqkeWKXLOkqrcwavx3gVT6wp
3v4wci5EeGjcx5QWN7jb6mRI+/ili3mGX1lNkQBsz5+xd7bhoeqQPWMpJHhymwX7EdkaKChxIFTE
VJvoWmS93cS4w3SPZf9etHLowjMMGcZThp2JNONNPT0X54ecsBI7uVrv50LFJf+AtHBsd7NYW9bH
ovmCg8UAZ2IvFZAeND4MfkpPYDDr6ovGAMHSzDWb4qn8T9Q2FZg1eiMUYwRlOyOTZmYEQQYiGB9A
n/eJCGoyb9/zGrqAJ/V9/hNjWhtgGcBAnGd2Hhi2yhyRfyBA7tHY7mk4OZ32aJLTSub5Z0sfQabX
0Xt0fG0rbWcdxRNv20+P/+1XSWjQLTlqoHUYZP/3X1xi/KyUx8bHot20X6l3+a4xrHW2C55XNYmN
/f61/m9VDRxuaGuZ//B+wluJfRQcAL0TtV0pCLgDHc8N9jdCFi4tbQlX1wCnUqcBLLMliE69tOzH
F+qLt87wSoBNKCrtWssY2yN3Q4W1dEyUKO0lFbD7nyI03qUGL+adCZdqYfNQgY4Xu75j6L/ZmuY9
SLgWq7rsXFP9ISeIKxx6D8CAlhpNwSbhZfC6AaCcCU0S21VxGYYwVLlPs8AuzoCRHlHWhCyyromI
poLZh9Ob2EWXGfIyr3vtwBh1SbcNcpfk5eWa5gLuoZuKSU2X/hvLRP8/zm46L00gfVZm30qz8Q6W
bdmwK0J0om4+ONiRFJ9M6Pz8FJh0sXz3CpZDw44gNxtG35A+bWNgyX/oHAbmdaZJI0Q8t2mdBsFH
JTkmr+u9Lv6w/ALBVUBpYcVZUmChrs1RLvbKpDO56D6Dx1jK1Ywz7Yj9wQAognK7yUCkPz+aJdNN
E/FZumtYf9PcoLTu5GdcbliA4SgsH4FO+kLse30i71vKChu5QoJIvCMR1QfF8joeHGlaDhLTZWBv
Bsowp9HzHC8fYYn/4mrTI+Z6co2rJZDcJIU8irVSnHE7v0eTeAYI6zccukF3Nr4qgtTfsmndbO76
gwwj3Vam/8fLJVPa6U/g7QC3q+Xu2v8f1trDdsOXhxi/iWTP/qbmzkQ9Hgpou+Ial0wMHi9Q9bq9
gjp2NufGfk3ULLn2w6QcrZnF4bXsu7ZRkxNyG7PEjuHios3Lz7te6EJpn06oJ8gSENE3kVbU1ODT
W0q9MHnL1KAyvglWlAs5dPXg1M6u+H/503lMfvWPesMewFAnpapCDnfmXD68O86TuD2WyX/nGWpf
DUIIAA/O0WmCpxy787f6lVCcs8GyvfuTgi2LAzVR1Im/XIKBGFlkSyYG7ZcTpkY4RF1gouWlYdF0
rD9JbzKDf4WEACt1ihpr73G1mGq4ml0ETpSvzxNzXTtK8jlUZsYcyIpMsmY8+rBGjqitGT5ituM1
Y5c3tJXP9sjkgCeGSVjicaPxmM4zGCsgabsCP99wJmL00dKkUM6mbcmUXPWYt4WVxNAz6iGt20M5
rTpZruU1/+Pz6591W4OZupjyvEkahx0KImrgNYduIK7PkzQ0WlDsPXvXGYFgMSb0MTqu2V4unHxx
9Z9W38YlLHeoNf0EwbD2Qptq1aAgoArqDEfBD0/M0se3LlZPfObIS3kqid5y++O7uCKttVqy31Sf
vSQHWz5lAt/yDDrMyeDsuxzEOpSkO3aVmJa09lZ+5jeodU5T4/SanxaYpUa2PnpJcAe9hhk2kNSC
nDDyUmn+eQ1/XGIm3v2UCXurXnF22jd1XgzhRCFPWvrzgPzrEwxS+mVQR0DVBKiEhmixmelrxL8T
+qOlUHMnIcFPeki+RMKxt+8kzkPSRDVf6VpgwSnT/SV9diiNTKSFSyn73LDywjTFuZYqhqZ2/GoY
BbeXGWWdp0C7kiIbtFag+DvfrOIQ+JhqBHQQXhiRKGK8sn5MZqe19Y4g917XYsB/78fpH20l6Dkg
kYgER61A6bWEELkCA1ecNJCWhtB6bWnf1yZkHF8Gn8+nBD8OBzFDZO+ar++IiBoxCWZlJmBH57B7
6dPGx6xysyWxs+LAyHB7L1bAUVUUJ7yBkrgDUFDYKWFbiE1Zxcq6i6XEY0/9a/AWBFjCQDAJczgS
gHg86MZ8L89c85ee9hp++P5ctpw2PzW6tRKlsRJO+nxcZukiFR45YzXkZTxKdEhTHC1C+3vwJg8N
NY7et6esagBks9zsgXt9Pk3cZ+4t2eratKFVZNt+Eeo5onHxpaoA8yscpLy4F6saoy0eb7K7c+d8
BrEcy0C99o+pmfSDeLc0SeqpYKaT7Y7GNEfEV8zN5y3Rm2Qgj4N/y2Zr4flTeyxDpaXGUOvM9hbj
A8e8CEGast828xG80Pk+dbiK2vAp9bgkQ8ulSJhueb4Y5pxCyhceFwDZpx4VsBG0036G5K3OhJT2
1XhYsc385CzI228Qi3nuFwuztyQi4VsZsaU1ZfgN/S1Vgt8uhsegGu8ryiRkul46t7AgroQCl1Ox
Y6D1ul0gu7GDw6O4bN1Gyj1d7uVcXRrZScAZQElhT/GOU4EJzTlrjfpbYXIyKJBQztG+TxqJYIHK
Fw0ZY4CyuKmfGtCtO2LZ4qkJzNbiXbcpAqs2Hm6icoOG8E+zwK2FEsugaOnOHuKcELueQOAGCcH+
cV6DNVTKLwcY+dwWYxo+PmNwFH0gV0IUft85+2/oyf3+qwk3JIl0jNkaGhs9ydoVZhAJhFfxGvJt
zvgsXrc2nVgQHfxe32jAebh0VhkJ25PfsvhupqC/knuGndgJEVsQSKr+BQMiMg1ec7iG8BiT4tgf
XSg9aoVTIE/K0tUcLmyVcfyaM0TZoEIitFZ31EOCVxaHbd3pu/BtyH9teCJjMN9DFDffef3alYdg
Y8JGd+UNB839/u07v1asxl6zJyzas0dLjcWizMrBG9UJ9Odx+5S5NAgUJUcWeW2bjtHucb93FvDH
lP+GYhAtzwQyJiKZ4+18oKILW/1OfAy+/ge1xCmrAIdFi2Ry3y3odWd02fgymK2XPBklAsgh8Kuc
M8D8t7RhaKsaFxW+SxL51nh0ck3G0ByZQaTNZ0yazd7qfloe2mFYX2dkpYbJED6OHKyfYiLjJNs0
/2neGXTob/DXFYLxr1UathMPvcZltJz/tUzTPz81cebhCfsq3mDD0JnIQ901SdHVMKmIg8qvErJ/
SOJ491n6aYewMe+0xzRCdJDjP8dbgIFTBXg5Uswn6Rz34mRofGb6Y95aRrG3DG9nrf4rQGTUJsWp
rNtutUWdcKpF7TnojhdeqwJhpkEVZBClTT5kfZjH1ibELMzooPCTkxSqSIYh8AiEwisYNQIQ0/LK
ljw1DzgUuJ+O9ZsnPTwR2fv1RRIDdgTU0EPdy/Y9mh2oA2yRQTPxUbHZkO9g8YuUg75K2H7rxrQX
yXoDhsUASWv13yu0QtWfvkWzFXYky4NH1vIHCDH7stjBAAuYfffdz9VuUPrI83hD8G/fNhnbOHiQ
/vywa/aGhVwqC636kDRpjNJuhuwLgez7iM5WrpD5RyJw5Nyw6U2xRbRbBLi/qGyts4t/5kGRads2
kvXReZyDRxNKenfYhtmra9uG2TEnNioSMTXOosy+HrlW1EDg6hOeOACG6JHA+qi9cFgzEyUdTXqU
0QqZrMaRJaXhM1Yob0DpZY4jNUUWkyx77A//oq4gnOc2Ok2cU9nopmM73RXS6HOFJtS0q079FjXF
6+mLByBmX1r1XTcwOuPOLEPso77d9uTX+6nV5lUfPFkrjYLohwK6XNLxMvop51kmTda8xFBn2zhp
445RxaS2csSjY2Py21DSDh97zVkUzIbl7aFdhnt7PPne/HT4OBGR8W4B4p87SGH4tVxRrPxNUr0b
JUHGyXTaS7qVRhs4js/FNWTgLWLbCl6KWwc9go5V+tWCABd2KCDT4vDcyAdXtXVlBq+vFcPfQtkh
scUa8M+Vj2ssKXqelyt6ARycSR/yV/FHaYN7AZ2xBMo3cvdL7tMVw5WhTf5vcEdNLcJh8k9KYkJT
X0ccFgePVGsSBVhBV3XoYbkmrlkMr3OH9tvHuSWmE6gc5W5dUcyhDFJahdbaQNFfAVW4slMbQ0iY
+pje8beFT5ysSNkQhCNTwekwrljxg8YpFPs0kHhmowa6jk0dVbE+LH+fucKLKmCtnfdwatwQ0wS0
In7jOc7q0Z/tbjEC6FCifUz6MBArhaCl5mMw2X/0q93fdoIZG8AxN1R6eHr7Na+wThd9zFveQCG9
w5MC43ZMtYutHBkT3BjjDnv+IeAXRGHASUajOuWaQeo8H3WJIWFZGuQ3B1yStvFadKSyTQkzgoFc
eS0ZXk0wv6vFv7wJRslTqMQa9beclhWgKI5fqx7ahSktCWduUZNm5k2Zl5aFn6BuBflUMDlKc9hB
04MMgCvNQx7JlNAxLHGGt0DNX5gyXTl010a0gGKov5WnI5D26aiTzhDcyuWjaCA2N548sje9zNCQ
90dgMq25wJjHKAqIGBlBVZ8jUtMgUajjtAnCQDSnNMXyhWz/eWRqhuDQLkMuP2M40J9Xd8vNfoFG
RhPg1CLe9A3AQuHj/elJOLAulfjJj4Dvhqi41MkxpzmQH/6oHn9dUCfmhyGuFEO7ljLw3jDvg0Gf
rAHBfK/ZHHOTpIfJ8WLh+9YTs7AqyXyw4BxNVc2XwWOnFVS068Eeq8iYOyoN4eDLteKHH02tmAwu
EACAoDD14YuMQXzb/PTECeqr9jY4HPDG3wx2HM5BzCxhLZAMcrllDgGHA/JmWDDoEYaNILAyEswb
VppQgWdNjC8clEICBzn70/CFH4Dm2bvsvWbmFFiCsQEaZwzG2gzU08DC3qwu+KqBCgbfSi9bbTfU
YecE7Ji8Id43M6giWv+thYVP4e9nC3Xy+RK5da46uxmbKinJkg7dEXHSHkeTeKUnVqcVsuBVezuO
mkHJ4oUl6O+dhPmVmjsf006KXUF4YN197LM4EGKzUFHsppX3u0dyJJlZhXPk8X0uqSgIupO6qit5
F0JBT6QLYooSK619G0BMY/O/8BiPtMEwSHaMpZ9SMQPZ3FtyOie/rpylmUGP/0o3fZBbMxTodOPy
FyEuE+UI7EZwTRBUgQoBGoSZgTSt6fkHpNreRmcOVN17PEUDwkKm+esg1Uza40cZH/URLB4uC1bJ
Y/dsKn/P/gd0b/Y0IcuMMK5J5WPTnwlfNf36+QnZOZO005NQluq4Ryt/9NFodO6AiBzfDUBqVI0P
jjF4n8uc4vtvvmW2FFLRLuEz/41hehaxpocmtLmdZiRbDUdMKA5+4WZ0Wn+WGZjErMPQqI4qOV/z
acu4btRXGJkrgWkh8M8W5ly9/7lScyrwmTSxhVh3V7sGyWsyBsPJxPetHR1q13ZY19nOfWp0w3hp
zkJykug1RzniJ67OrckJBWbrHsSzZ3jypQeDfsXkVvdAYOWEeBzP45NGJCfZzCocMsaft+A3jA9O
lH/hTHEorF2U3UYW9nC8zisr9yiSxIsl6sKR4Ew+h11psakd6daPCRmULWLMbxHNARN3d1n7ZrBQ
0CJkajOTSCnzcChIEFwt3fQydPvcZ8ZxePYhjsMbxRQSS9iqE+L6WAD3d8XqLw2r/UaatHUmy56Z
zWZeXpj11l2Bcvdzb/PoS3uEP/74ImdROVc1jZf++qPwlAO/D+1FySe+643I+r8fxlEbN+drIkln
wMVWQasnMGP5yyXePdypLh7EyWVxyxRFjdPz2FWtG+RmmqOHVRBtRRfzA+aD1q5fMZiKawCGZ4UK
kKmfTfw7jhze21eTXAVIubb97SQBagsTUIznyWuyXdq5rnlfUV4bwGVb7iGNDFtup4do99WJeUGO
3p64h2N3oQnzvgLMInjcwdOW3sMZSAwHuG11omODGVEiYxUa8HynTMRooVghEuPhvYywgBnA6mEo
lCEvpov7TQRXrRg6mfiy0LWD5YLaYlZXHkJ7mGlZM+uW3Yu9hDXOgzg0u4ELKEZrKfreFUiT2fJV
ezdwS1xn5vOrn1u/nhT2a9eLo9WTL+PRisPoqK+GDGtIbcFedzmeWbZKTWvnwjqA74X8pDPepd2R
+m3PPIlYsUH97YN5Ke4q0int2QdDySH+9MnWid+BCmbzaqg3TSOVIFzIToTG3anXeK8KXnrxiI+x
Bi12J47ni+MSAoV8mPo5zjREfaMeQLt7JECneBTFR1RjZgb/vCA9PpGRh9JfNEv1KmhDgsxbB1/q
dPS7W+G+78vgZwyjVAlp8GX0cpdOUJ3xJfUDWv8uZwKec/eqRO0Z1BdKJWRxgH6GJany3Y1Lekng
jiK4FCToVQjzxompwXvMKKeYe5RplD49+t+gbOLuOXgOhFZWr8HLMLD5Ugt8/pQKfdMOoLCj1G80
BNnLft4PxwKYEKMePMbdLWItYKa68kYm6DLV0+hUaeE8JjOtGt55Ku4znsoFB1tX2jv2azA+xqXQ
XvLNPe/vB4CRCVUeM/nNl9NC1Z4eFqdq+sEm9ak2jhuNSfkvME5xJpK+fcbBYAW9HhBkcSrZaNCz
UzRUXnp2MRWOFVzq5HiApTJItc5vXTsfZBZaOtCfojdb0kyG3gyWgP6THZL/Zun96IbEq17Gkgff
nrcQYAuFix2gXzkGPdNaXV7pZoJ46OQAWwumuRkjD9uu+mtublvw9VmpZ60l3pceogKdIRto1DFD
kvkMJsG1ddHV1O0TWhBkNPHg39Z8OWRSlqwv7EFWqc2UYv8tZHpoeAwSbEWZiQDkc3JKrFJpmSLK
yXAxvk5I9aQK18dqpKtlKqrvSUMijQLbm3WBGt5e/9zKCFL/cnSAFrIN8R5YC2cL9wlGZ3K0xwAV
kP5UM+XuqEwyjn5WoMsLYvHtOgj26FW1nlzHUMjP9YuuRpt4dEYWNvzas1HtL1OUD5W7trM4zRiP
F5mK1RK+LfZzhSxDhNmQqHJ1KveTk0dsqXBckVQNEC7QeQUXIM3EqoZWDlJuDw8DpUXroLFb0a2h
NpEcGRUni+WzacfDHMZbDoOjia5zyZ8gP3KaFMdvzUjvBj8vQrY+nIAZCyHyrmFcgDK1JNPMzwWq
iXz2rM8+gvGOfV4HAqwl+pE1YOhQNeEfPAcvo27A/p98cmQOziq8Rk7vp2t6DxFzh0D24VuVltmb
piDZB3I3BEgXLvKgnDsPLmpoUqrW8Rt/MYRmk//vVRuF6YEJB/aE66Dxol0rJ11v1sK0WO1RmgSl
YT+vZrhdHE0D4BW3jur3x22/lF1SRrJYWFIrEj0rww5YtF5vVQ16T8WC5lGQrhzoxRpGLMLLlaSj
gB2BjTekUurnkTJkXtzYDeYHPRnP5lwnNNOD0kBBuqIq0ioL0cp46MwGzhE4fk93df/sZNXEw2z9
fwtBS4ZiH9KImdAJxTnjPDziz+B9fcDA0GeDhujRkW45V8SgpVAv9zXpCdeDCLwJ/7GwtzufKVBa
Vab5ywnb/MxwCOn6zbzhbTgdPMVzwxN3PSuwji4bJ56PpHcBW96tKrlam7v51OJgGAu5p30I2aso
L0D9FbmkOuNagfTOyWji2FphNmIpvvvyXbI3WULeJ3y0eDalrIGvLXEuxr3taCThpsJ5jBi2lWJJ
GNau7kPLv5TuEzSiKtkpx29dYUr4Ln3YoU344NT/xTlElttdWeKj0glMlLLl6adoeuHNuOpfrKB9
1o2SLZtltzLI6883DkrSNZxO/NFi3WNVbxgKU6W+B2Kc2KHB5g5TtjmmFRPN1SwwQpaTB5aG6gAa
wtNkOnatZqVCWjKpbqaVxIrSmSElxLxS2+DUI7FSEJ0Q0rEC8Z2/qRNidBSwv2cRpjZZUTYPbVyh
8FqopzjydwV35NwqxkAT4UtG2cAzPgGZUwHQE5dA80w2HHzxF2qDq/2+2yg139mjMoyaviirYJxp
jL4xiBa6m9RKsfoHAi8UB7FSzjpZgpOZ6jXgk6aVacX0W2JrSFyYXq5O/ZP0YZSu/XBTyY21avUF
9Z8JD2TMtmTN+yWJtav3WLABgpYiLLbLVSPbCGrKeFPPtOA9whkkgP7uTEHGjmmsyuIR+FtnmAsz
bQ6sZ+6Nj0pULu+ZB9w3/qnI9uR/1iOrVMaXlWaIKMyP3iAavzN6wRBwIoK4GDNIAHMDEIG6T4DI
ANFrCP5EvcAKThOwOeTAHJi+z+d6UKCs6KsP+awpq2c0TQf2korLNstlUPFrxQBJ9/m+ZAMQ12ma
LXgcscmnMqfy0a8iWTa8s9sIISdgNaHlEDKtlXzbXsacqb+QrNwu5X/C/HkgyNA1H8YcunD+ckcd
9Yc+i99q3rE/59YLJ9SB1QtAODGwevkTGfd/b6NNiVeHkmPjSX4I6ir1DuC2SsEyMysGaJQw205q
HeYEt4fF562v64JHCQfpPasZ7XmpY8I2LBigj9T6ZqSZztD+6ynezamfAvM9piTES7yTYM6aLAC8
9HVez9PYV185DPwlBFgTjLV7OPgXnN/vm5BxXr/MF+Zfoyh8a7ecsLl9NrfHfEoz1cY2HeNR2rmo
BCzqsA6ETWvi7maJAxKLtIcouif7U+xzfUGFCR4Z4kEocLsDmFWwX6ByLxrDy4jPtpfgM1ZPduPK
kODsL9bhTtbhhkQS9u0TNPAj7OjcqiMX3r4HD2u054p10HxBdhyxiXQnwXrnO7rDAYcmmGOHUpni
xF9SCRUS6PIxpXjS4zUTQ9odjmXKCXJGAyM+gFSGY9RWacC/x8A5/maQyG2MyRpnBCZ5nJxZLzz9
c2ea15c5D6gYYnHITgRhaXahGZ0uyCmTA4LzC/tZicRJ5FVbVBXDdR89S0KshFjaxa7qbmSeLjW0
TwM71HKQFZaEefpyzU7EPggdmsj6QJFdeC9CdoKuN7N7D+w7dqBwX/SZgry6zombSU0pSWE4I4Uv
U0l9/JFCNihOJr2HaA1WiY/I48f+THyDYIyNOw4CbadhLeS5YXVVA5akYHKVDP/hO/OYhiMOkhcV
nwKfuWjyw91eSGpH/CEdcktcpFMtKrusrXXR2qY5WfGA/DMaQPm2ViQlBp52vC7aHS4GScLums87
yB4iYc8OFT6PyJ4XnbvH3TQHE2zYZqRtxfn6hddcSdVDV/3OQFKQ/o6Ke4xe9/ajv88mtTJXEB2y
Mqbgj0uJhJSRPaLMmmLWNzeXDpktxWFm7VCH17fpmvDVjYpcX7YkuiPM32HtlWkR53YuJXv29QEW
hK8GVc3YVX2Rkz1fV9/SJIWRDipUghtXvcydhMwoz7lFoGeoEcf1r/JKXj4DWXSYw9V53+0sFiN1
Yn6JT/gLexpD1Idmtt4DIQKyxlnEYKoStJGC9UL/bP/fjIuRKDz6MkAFD9IeJypYd/qSDirPdVSR
XK/qJxEKDM2OaDwvB9BpRxWHTXvl5B9kYt5pT2DYPBta6PdiyozlxcScU1GAR74vK3+JkSaR/1d9
O60uygbGzlKG6NNM4VFnlZttg8nCLk0NA4xGX07yDI5WeM4eUleVos5tu7jQDqpBA4YsPPTUE/NI
F5/ug0ujdLDFcgt+DQ4Jza5FEhmiWhWWwmgtW4p8rsRPJnxXxgQ5CSgupcT+oL1FfI1T2xDbB0L9
0d+m6fMHhjCZ68qzmKwyto54hyIwusoqn34wdVdc4bbbb5qa8wGmGVmmt1qmDeWPKVIg00skbdSz
HatmHDp3FDYBWzmPSIjOh4EYnHdCqn5Oso02DndwH1T8SOVQH7QUIPS23jHBPad+97B5RhFfhXXa
Au4N6G1fM8jBrlk5Zpv8wHUsQdhbtTnNoSDDV+EeB/3kPzMBoRW1qrTxNNcUg9bvG/jA+m8dgMgh
8SJjz9wm97olKyH/LwmBzmGLsT1Z+GAJlTrkc89yPaKQ1cu0DxnvX2QsVj3i30vSy11qir3gcN1R
Utn9vBG5bchMeVuBSVvClXs9zUGJA08IsiXiKnI1JYa6v/rYFQ40hXmlzehbajHmKgdFHAIwLQyQ
2O2v8ppVElXAIMxFWTZISWKm/Wux/cidb+zuZQQEseSdNKf1wpFR5xzgile1++axNkWPjuN57gW8
Drl9gZCl31D5Zc98wX4as34NDCOoHDiIZC0OqcgUL+LRYP7SLVHjNa+xeEmBF9/TfxHlKaihBLtz
gzWlEGXy3nN9yuDnENz/FMeCeIzycFOXvTryDbgxzFjTfobyLaO0iduW0VyYhnRDA9dLHfZbz5Q6
ff5LxbW8Ia5SHLQLXY6s8WHRrAdGRttvRtPnF+4eAueqdZwoELzmxTDK+kmnsuiRgbxjqOZOsWSo
VxH1zBanqmBt/hbbdAL1WqihR7k1nFlshSCijNTUyvnjgePw0QfqTKO5y/28RNy2ZH+icEviKFd2
XEesvgxisoX68eKXcgIPGAfaujXEFUZwnhRo5uMs6qnDwmaGIFLxDRVCZwR3mVhAF3DpZm5qrxVl
nqD/StvMRadURZRLGPIIvRENjx3xlXVUnCKAJjEQ+jEYEk7hBvhHbPaBxaLe991qW9FUUR/j0Pzn
wzEcefPePjer2Qi2cARLwIh8AFdHYCWbABchNCeipfFM2TpqUWm43A1gKdAt7tzc5A4FY/oMl+T9
J45W6bdeied9vIeYuaYpfVnLezhqC+pt10QtD6GE+hH+BzpZYp5Wq7ncLAk5UngzGpNiJ9/7ceXO
e0AuU2KrBerTbzOoQn3A23G/4lfFVEKnJR7N05A9jxoODWe0XIabrH6UvukjVhu1NbG0SUSvGUCF
cpQ9jhPQWoeNh9+17m6ITjmXPXqY2JaJfPmtTuWMgqW7xaOt0QxYOjOtJxKm1beTqOOA0oYAxhAE
D/tC1xWm0QzHngpIwHZS6RvGDrssQoSbsrMC/AQSgHi6pGdkvnzVl2EqSdWOahCSNkAw0UwebFzE
Wdgk0Ff8vuWGCr82xQ20maCgNPeTx/cPJyZls6yRgQx2SWwtAgUdH4qODqDSYvzi4mvWllMi9iHE
fS6UbJJfql38HPIzxHIXOfYtFMPyVWXA/HTnpC8CBGqTcKZDW/vlKV6HIciTloDy7hpiJwIN0g/a
7+yTPewgWx6IF/jJz7SN0uPaBNcMvyPJisNJc3XYR2xvxKb0NtfjkTiyRUJULERg+R3YJKHlVfj+
WXT3ZId2yixO9exJDol3KRCyOThVJtGEP01WoUS0arD4G94UMKmwGJNm792XDzu2INmiYT0tdua+
EU2cOEaYwQ0eO2NgUc8GSIaoYuT4l1ULYm/3XtQze1Aal/JSB+YzCDyZiS2A4cuir3mBKnDz1vO8
tj6UU9Wie6nuU5oBLyqTauwqLeHsavUxH+ECqdQ3BeQtiDwfezbi4kKG5zg1G+lDDS2TGlTYU+fs
CBmaMInt8H71APM4wMRWgwzVYALroAh5UUTiR8AaqLldUDmBlumH2idU+03E5csWxnwiOA08kKoG
GTqENVGPUi7AbBOv8eM8lAgoWdWYmW03h+Fr+FW5I1Wk2vW7C8OCOuZdrH6q/OskmQOvCSzVe+YQ
uflnJ2hvK47fAQLCFpZoEC9PZ1bVGnf74cdFV4RTaFD2IwrWtkNykVmietPSq8R1/9WgjZNU+IkN
vfWhXf9mn06A5kfai7AJUgVNMpMQfefWL1ZqojZKlbD7lADq9qFYYnWOEF5Y1h8SmN2yBPfFyp6Q
dDDxBn4KX5LOiFWol7VxrHcMCKADKgrAV7erD3QTYijULjkso0dS3pgdSC2IfpkvHVmVtc/siUyn
/CKUN90rs0am0CRjW1ms/QFIwyHM8JWeXOEgZxFE7SUcQYIbluMoc265ecyT7A6wmme/QH+jeQnm
8wW9pWCWgO3wwpQDXfRIw1DX1rNpNxrs0WgV/glG7dEForYbsIrJZ3g6jOm9J8xSJzGs5xXbXLmT
8F1PF5kKF+kO/hmFUVs5+C+sEmUg+yEunjVXdZy80AV3ndxX8VsUiIlEk8VzAtLKz7k8W0YpJLaY
6mfd3vJcytoziN0B2+5IlyeoHE/ykZmlG8j8pCOQ8ONwlcL+y/HcAI4zXIR6mskiSbJcHWAQsSHY
9beHttbOq7vvNfAWV+JPFbEBZ9icHmKMl2y4dwG/AucZK5Uu9BLkpgaFV3oqhlPSVNqMexCz45JN
9+6LqfHIsBdDrSQ7wEl6LFGq8ZZ138g4uBAS+AJ8w1koiZz+Dn7GrCFp+7d3dyN+yW1J0L7hoTkt
6rfzzBgMT/vbBL4v+zxX+S/eFzzRGePkOXzOzl46ZszNysZtN0VsBrvJjdeboO5qqxlbePf+gl6s
1a1N6FpOgqFduljc0m1rCIxWlGBAb0CyxAkzQuptkoMFr7AEamx7xJQeIDZusmIFgBP33Lb6SVo5
0ByvApwPyQXobz6XH28wup6gF7k6y/TEmIzWp5jubi8fgiOw7dksg9jZaLMGwUr+Prn5wAeobrho
pt51+rQKXIIKKHlYPtNQ06XquA7/ALmllSaptg1lm5d7SHJb6ZMJSR7oEYvb7lo+AFBjPF55Yx6g
ffg4kh82xubp0kQcV7y8Nj2NXwqovCOHaH4JEKecK1dIfq+dZ/IlIEZqAL64nz9iNboBpJsjSJYy
0VQkIaekP8gd8DZlMKrzhEF1FPQ4SzzGianoC0R2KC7GZrDpHhaV4dYvKasBGI8Hj+6zMZROyWyU
lD2BofzgP59gbpJoJXV+MkyulwpWpFE0/m9AdbZ3/X5hp4G5TFIdiMZhYzPRspquyeXusYrk/AAS
U2OAb1q9wRe1T0spWutA392MbK1iCb4ypCliL94pzUTTis+Kv+3eS09SxF2iB5UNp5u8Z5vR2ZsV
2pWd/louJPByVYZifbsyi9w2lq+BNvk6xe43gnG3PeufRWBWj86EW/EiGp4QeqtOoSre++GXZEcd
690HxUTtCHZv4nE4S7xUa5WfJw4uOo1zZaApew1TnGXOjnKYSRjwfYCD7BvwVnu+tTezZ+jeRYwz
e962Cj13h9vU2Ip6OfZwRotvp8SDqkgoc9gisq+Gb88eiV3B4N3+BTmoKU0pzlSTWkEj033LTA1s
HJg+fjp/611jGMilvLw4Q9Qcw8+1roQwUalt54zu3psN2ttrKWX4U58Gb7k//V5pjhfC/3Cmi2r1
w+qxvXCrIMvgS8UeEnFphkAn9RUzaF0Ywk02zr5qjXQSg+2qa1+3+x61G14fQxj4e9pBWpxNeeeK
b1Q+jfSOUrv3xGFxgQ6tAlI7Ivipz0/72K8agmw+9HZjzVu5mHRyDms9DA2VtbUj7op7o8UnmgZX
27cfSdvaW4CdsMDMUP7zyKzTNyh5w8NN3ekSdnbFDdB2A25bP/6wA7JyU2Ayo2LSPHd4iU5Fp68Q
EWdmxlGqOAOq7LHfOv6mi1X8hbPdWSvRYgsqO4KkbVDPci9r2pxatrR9bgAeW0qyBgweSLp51LGV
wkzyRHA67E3npk/ZriCykOg5ceiHhGnDPM6LpWrXFejToS4r4eYlAHoODRMn0vsTA/JqiGrTfwNi
VUqUSB/IArYLyAfIWDGnSUwpumlVt5PaBEkk27LzfRdb2Sbp7Lb9mQNYkvpr/1SndSXibRAcpznS
1kSOvojVPBo6CuIuxc9iLYq9lWl4a2VKqn70i4EOunmj6F5Oyge4zsxcyyidw9Dwo2nU64MNIY9o
qBDKh5hNDIKN4XEIUoMFflgA8FGFlwulcVeTKadf4tattqeVsCROViiogRMq+w+f1tzoAiPFQkA8
ZeUGEhPVE8yPpOtKMksSjLIY36dm+39PcEtDkL6ZC+8mMIrWw+0ZueTWO712L2RZxqnt5Gvsb9jq
+4pC+TBnicY6YeQ0rJ9oiwRIK9eMoPsEOcDe5YaQon8wELsEzl0fLQK3t/wDQJCxYMLKeVW5fd35
XT9MDViIRTickOvUd52y5KVFwvEkRCwHCDHx7aGiIa/q6fyGZ4GMD21GPUur7JZpjtxNsK8PKM1X
g0u9dIDW45KfYa4Jvjff+8wMj0dJycUOg0gA2WtmZAUitlyTHYWsL/ulxwu/mj0Jpg8NWlm8bwdt
qj5K/bowFzZYuCu9scQRcmmsL6SFBHhU8RsY5KOig+tWmeNzjYESSMKpQQLU3FxoXWW3jq9v98pM
MsJvyBCnV/aTl1q64X78AwcX4fW/e3gx3DY48/whIzq+wX8Qo/3rFcPmC8rz502n0yHz1lzN7kQO
xGTboFnPXyROX+yit/0KwpXPovoy4LAqiGDNGBzdOQUStcbMEBuz2c7j/y5zJbRN0YLH3L3pGPfj
Pp+ccOidyeNQIlXMFSk+xtzNicl/jtf0RFIeH+dEi/avc+m+BYQwMJmgWC28ILzHsHxaMfwO8y4t
zuDiK4QEsvFvuHFBUsJi0irUU2x81uv5ipmc4U6xLDm8WoXRQyhd/rG9djXsuHuZzVGGg/wuCSHj
9XFF3VblWs1RDhwBsdWA0XPxsCK91ZDVN13P0KJKsRRbSyMfOY/HZCQjWWdiaE68KKimPGtgXDVr
dm8OEnOTHK7r1RM874a2CkkCz1dLdjRjJSc6uqMwyvbRMUMaEtpzqS0psOXs3mLHL860vK+TB26p
biFx+b0bRciMTkAchSa98G1Cvi6RU8H6XWMndq+PeSxsaoQj3+KxW0S+8USK2jH3k80jobpw6Rr7
aNYaeQLPUM+q+2+VCJvtP0qOCfQvMHMfvkj+ELbf3vdtYWu+fafhrp219r+CVeXfjS0oNsCxqQtW
7Ps/aWLYUzgAWGC0AojEk3NimRIwEbQ7ZYWbzPFZW2pnQjq9aP4kyWWepA8Fx0XahoNNqHA88fqx
v9eR0ty1Y0ZhRRDUHOuw2eXm3ci+VKeuOMivEEqes+AgOvT7qH6YLY0zf25dYk20+bYvn6WbLKdN
YvbpdN6Y8C2RObTzRlRjBR/aSbqTYXBi1FFqvG9pbTD+Dl1yzpZAI60//MFqYJFplP+9rW6wtmBt
25qGueVVPBLz1tzMbsn2QgNgkeiOn9MQI0dppumleEOWiRghapuiwGZZmp4ye1YZDOpfZMg9bDpA
w1Hjo6Pxpk7LDwnf+1ehe/ooPA12mUUmRz89a812Jo3P7xENSqMBJKAVVa2nXyJQ9TYvWS8RMV8L
YEtulYMoatYHrpI9I7Y1AcXxO5ssBpw8NxLUgg9d34tEyBBDDHMAbEr8SO1pKhaP0MdRAX4cmk2A
wWnonAz8APhvYbSmmWW0OCWRjP2uCDxqYoB4L/G0hXCinZ2KoPXQPyITeehSkAnpKdm7SFSf/Epa
tozkmti/cGv/q083yOjy+V+VQQA75E9PwppOj7jsv2KmQSdC7mHlDpn2GocrjgYrOA3Az7VoHqcQ
zQX/NNqdAmfrZ4ZIF7oxwdVQJG0ZObQyGHQ1iaYAuQHBcqP1MgUOnPNdw9Db6ooTl5jMXjwbMQV+
trkbeEkEELhsI7SaK8V67V9x2x1MTLDeemUELz0SuHDdQnRBxqOYNDky2LASoKnEps3rNLBJgQfM
3O71hoooPdK7RF4k7CbIozL/V2Caw+bwitbOzTOHckhvYJ1yaqa4AsWSnhkRHjV5d4S+JLNem55H
1Ja/pGvb9OTkyiOhzapEF4yE060B2It/q2InTnoLHJJgOIn3srhP2tbyam7O9nw0lgiM9bYIiZiP
4qpbrpoYFI/XQbHXR0dDsFHYhiBUDh72ygIHB7v9wPmUBYBConulDyuexQ7LB6kiyJX3FNc9TKR9
Qk/YEvWYmHr06hdwijLHXM5tAxsZC1M1MYZNqPYPgDENM9QCELeSSMOkoN+RcN68mftvUVw9l9jC
E7NlPgvcmTDgnliNsH7gkLlKd/nr3yGw6zX9MbQ2abimW0Muk4X317HRKxTIpSwm8y+LijefaRcr
I5ASZjhQRfT+y0RVQC8+n/UMlLFY0UTsvMRc2O1t/3zfbJrHpTcgdA0CbHfCAtKu/5dH6UKNXLmD
wXtVtjIdHyUQUbz624yqQpopak3Hl12NRX1xYRU5KK8VPm1KlekpwZeYZiezw0Exu9IUX5j+96xB
BqboSHK8jKfKhyg9DPkhUQ4e8A3M0AFdzuC/15z88JEwaeKjPE1CC/ZeBk1FC5rLeLB1TlkZO/Tl
CnmSdASGPFOY3mz3nL+hDd/2TkiFQ2YWzwt2hB4cEHZV8tzabOjfcwAfCfkZpeQPKWK/uQ03wvJQ
EpJi7B0uQATBai3yV8WmGB+31NmYAl0c2WCtq4ypwCseLarRorPySaLp0NSs5R3acA98KnyYZrLs
K0PwmQ6FPeT5Vo7r0FJdjHGqHeravOIi72WeOxYQ4IDayRp9Aes+hYQ5YhC+PFAK8+EBepRvhv9V
6+8d2V6zw9upKUJ7tGwx0NOq8sFzrOlhTxaTxQHKPlXnV/BpST0ESO4iLf9uQM0CRGPvS1ifRsrl
9mDSs/hO5tMpKZ/ywnRmyLObPeYgaLrVO8QKoEGsWOsJHJ3EsuYySWNF4aRVU1MY3dEncwPMx3uz
Ktc9PhfmWXHjM3Jeb+VCMTD0GjdzCn+SC7cYMncyHFd+ES/UrI4Lc5WF1OeBNP2AglPCgewK1UQq
9hIFTqC5S+smPcaSp5ARfnsDaYgwxOdSBBctF6BYk5Eh4Z3v1XbNwcMXhaWVOaZYUlkc0sg8+fZ8
znF4QHCPWfKUB7w+TKAm6ae7qKj4t18HRf5ouJucUPIQ406WZ8syBpGGKSfiXBP91jU9do6K0ERU
PZfZUai8yN1dl3lkWEZoBMuihHmEsQm67n9GWqDaedsna2fyKtx6C7xNQZBQPyzrTXprzEIBuVZV
sE0pwBjblH1HxxfvPZunjP+Wnnxmn3AspgrIetLZP7Mb3ISY94NtrM/lOfb+0nhdC+iPbi3k4+j1
W1l3TO9KX33eYbqjVN5SLRq/mFcI7+p4sJ+zO+TIQHsv38pdOGt1X3J4g9e1QHGN5UpTQf5Vmnf9
GBZ+WW607ue+zD49sWPOra2vDXVqRS1M8VG8YSLfGzVIIYj77Go1hHPEyOl7JLTrfvTLra5z4hy4
AEP+YCsdqP4dyAo/cTmw4rUWE15pjZiS9R31v2TysYVjQ/+t/6GtVO0XzmR8PbSJBusKGNbEpwsQ
yXu8XjN+pPFai2vC01k0N+jXZQuE/v+cuWwdNzC7Z5JUDIrhHqasdt4+gbpzOxM113SW1Kn6iyNF
IkJmcXxw7KrT2Adyv5+ZKDqbCGNEUWfgn1KxpJZGjrMLrMuUsNqWPf6+KgUzAKOmV8dlmwsedY9I
oHUQg/AQtPMDwm9mdmJWjPYENGbQJZYVQQ6XOKAw8GfbuxNcP/7YXYolfpjbhO7NWWdSTYJbwC3A
aGRdty/oLGCbjY09UiFzamdGWUvkA0jDPPqgVXXCwmH8YNU68OPBQ9sIyYn3gN5lhBvF7WO6PhgM
tzWe42vF6SAdZO6vC3WOn6JYp0xzccF7Y2B1dvzi+i2igYOXLK0rmBH5+1gF1WcRcE7XxR/DWcnu
L//GSkY/FsCdTNLtzJ4JKvOcZTG7mpCbORodnuN3h86hntf/0qBzBYFtkdf3OD5SdwuD89fP0O8h
IceT6LWtvEwGfXUabsmCLiB8sl5R0NHb6DVV0WsvWmQmwfjZyQIDSYpTyxko9yv/SkZgY+l3qRNV
PHHnHG8ZL+VsQl5J0+uNf+1OCGzgFT/tki0/BBWMJa3Rrx7oGKmoO83j0e1DFVKUMbUJikFRCo68
hIvoYM98C89h6Y36fLhv0HVktEHbToCIJsRJZMDO80jLjFmHczvapBKz910Lfxzy1VABrojNXQqO
Dc3u2i1dI7TrvdUZt6XJpGDj3eUmRVemIXZODZEJp87bgzv7jCxm29dltOy5JVYeQ1Zzc8+5mg3X
Pww/TCfr+QSU+H2S5hRBatTDALuYFukC7exZBUtIgTbZaOsjvdtuOVdBAStBeBB3IQu0+Hytjnlz
MCHcO1PYtYFnTCsAYgXmGVK8eS3EdI4W+xJM7ExlUKN0RLDR/dToW/dra3jm7ve9OfgJG+dSPSkZ
Yt54hPZrGZwBzdsmZS0AM8eBN+M/BBVmnFpjiOv2Qu3M4OCU3H3N3D95dKiHgz3xwoTIey1GcE57
JrfR/BA20WSCSurb4xO5qaeShPyDRwEchY4BWF7Pcor/0d04zNEVgRfOGZmogvpjCMJEhZxAZiYv
urtvSvbWDnqkNMemxXzEgEZRNlnHSgPWa97bOY/h265bd3+/KgQc86wV7HOtTaJVzoC3UWWSN3Gg
gwzS5thT1slJbeIOhQUeHGt85tJnWLPnn5CgHrvWGVSlVya2VHXbZkvgJbPyaczscSJFKkLy5d2j
MJDosuEGJPFZ8OviOy1S9FVvBM/+38ug/jpwSNA3dqQcvEFK/GspWQG44zP/uwsY2k0QEAiUZM4U
TXcpj+uVuI/mqQzQhMJ2mWtfV2fVFxn6nVH4fK4YXGODoR5zB5j8MFkuiDpk/Nw3r6XVrwrSIaK4
Bkqj9hjU4Hfpx7Zqi57eAsA658l25fcVO3PCavh9SStNkP5oGlgaPfd8osaKnlCwbjLdVBHalT6e
YLkXMOm7FCCqKJtPLiSMecUchynuVlm4H5h4q1TRNSw6PkywXOZVLYeYD+TJIYyzIFDxbMMbuX2E
qV2aXbveLqQz66RWESV1JUOR1vgjecTerIkGfe48LPhuog5OS8kUU8oX+/lpHIOzXet/54mrVpcr
H06ipxl35Iyh1/xn8IJqtHSaDXHaBlhZ72jj6yerjPv2nNQYgQqIWkUE9asmXruBztRWacXXYiF2
P2QRLO7XbXiVGWN3eXfuPI8YCZ4Tf53KvlPtYzyiekBDQbcGnSoRFsx6GPraMpo4moP9o06dCZA/
FofVKJtnK2ZqLHAcJS08XyErzSjOG4TpU+I9AerGARCHyTW72U6OoZxkW7SjnRRkzus4/3fk9DKA
kc/cvG9GtK8/1bsVufaS3p00abEKMqMTg6P8xe/rXcWSRuFSB/FZN75Qy6ruT92yqfBrD8cphlnP
5xjdFth+4wm3om7zXr0v0+GvJYMUTE0JYGy5WPNbbHmAzFxBRf7D2VLAdVd4pTMZHrO2jzvuLWip
bs30KVlzk9CYej8Ful6CQrp82yPeM1XSzFS8f9WPSxqfzv3UeNcG7g6y46jdZwl30CQRh4iW65B1
EaVhN67TFDO6xFa/OvknbIR0arK0WpGVe4+0oA+6213g/D3L8tFKlYrcGxOuAQr2omhs4IF0zx0t
zXSiSO2eLYBioCZORIHVXcCMCeA/HwWNYD88p5MkEyUu+uxrxLNX+VprOsLOAYHnxQbCVJ2h0LKy
gR++wooBZtoND8zTHCYxLFXsXY81wlyNm2FxFxHxXyDn8yQolsPjpEFo6ork/r9sRHIN72Ffbax5
tYox26CTn8MKDUgp5HnbfdyuG0bRvG4NqJihNfZmEWdBarqgtM+n/CAQmEHlvh1f21M8LnN4EiB/
8hL5s6BfqlPonqixgfiHe027W1XvJk0Q8x8exrN8b+Pal2u28CxEW9xVuvkh6dMCSdTLAaKdHXzj
fYFbYm3jmAXqOsVPc7R8PkFVF8bB4r5+0bVJ6I9vVZ5ey+i7XfV/cVIcgLbeENnodyu9LNlXNc1q
JeiOv2Dz9PjWzOKeD91sahJ6p6jl77zpeHs6DkR+SYA5T4MoZFodZSb+C7VbsQPd1XLsr00jfkVG
4TRAHdlaytcGKFjmp1azttVWGgXYqzINCA2C3nzc7hnT6R1e67HdTdRSCgrLuRkw83/iSbNCoeQ9
1SgjuKkIKJUVGpqxU8EefPg4JZwjNi2EajxvOQK+ZTpkqYTU0yEy0FjApQWgjgd1HKey+HZfF1FF
vCYnvvxvkRyG7R4Wv3VqdviHimzX+D5maJshEbsa2OT/yEoxEclUGSmjvpNS95I66VcDocLE0nak
TUlRGMFuw6sPnJODId6a+u3PypYrhPq0KZzv1YHhQL06I6Zz6DFJuTbyu8DxqMUDbC37VmmRaxAf
0xSRGQ45nbmPQdp27SA6PPV1CAUju6km1xeM0u+D3k5eJPi2TrqgnJTWbwmO0vWe4zYhFL2BHZUC
H1osHdTN0JhzJy5lUtYo06CnwSnSUJwzUAfvo6AXu7izaZ+2MptQl9xDMm05h29M0jRyFz1Ew7v2
yl80xRpzVNhjgn7g3mzjw9GMgN8FJsbQBSK5yoit/CyH79dv0bD2enENof9d1zcDKXZUkY9AG1Nb
5YxICGKBXT5doeFhy5+GTx7lpaNp31BQvrgOKiOUWG6UEzuNxaRU/CT6EqdKrdXiLhcAt1cAjvlM
feSilwhFuDdjmJPlXupAl3jafDwWXZvSpAoc/9pgA9qsxAG7KUTeGFYm+Dfc18CH5dH8e9a9uzz1
yetZcH9GpgJrUPbUghlKIkn7UNmr5qdnwv+B+5t2kmQPRRV/f0vI66zgzQZxRzdPv7YzZY5iNFSY
yHFh65+QLXQT63+muxd+IPSiHIaH7B8Im/xMgLDmL7oX0vnX59XQPSindvC6xkoWEMIRgKrp/hP5
CPUaX/9wxb7Gw0no9SpGFaaTdNf7xge+3cdsjglvONHY9rQKiekE4MF/zglfH5VCjeGnuKrmaLhe
SxGa05bKIwmVi9suW8vuHqVtXgSnzRRAa1EoydQ9et/Hq0Oz6hYZyEe6LSTiedIaoOp3E6KgBoA3
/rtjsu0JUWzVpAzrvvrkdnx0LJBdYhq7k42Xm4onak47njg8Ku5HzZECk05ua3wwP9T3xEef9Kdc
C9bdCsg99SgKdni7cnOQNymIyw8Wu/PDoLsHxuoliuVaL+jOe2/96LVhcN0FdAfV9Fv1b3x283V3
X/PM4mILnKv/PcnGQCOjGJlnNm72gR5/OlG0tS0GmRSGjSYlhhHN8COdr66GBvvpCDsRHC7ASKOF
ok0k0wtGroraYvsWhLLkXx7tc04e0pFAUjJarRFHx3RyBD+AXip4VVl9anyDYcnqN9i0oOYvB1i4
k7y77yNHDqV7/83CsRSt4mHO9YgzJCYMiaVRmb3vPjqfY/ClFbbno6j03KKVYUiR6KXVhL/Jbf9K
Sl8bBlkVqsuT9UoH1ZYKX1iAyZwdRBOW/csZfdNStG/rMi+WeI3slGLFnjJQh3SLX4VfGWoGmr6G
yoVTofR3trLBIEr9RTyI8p0oERJ7MyIDxzHyxt9pW5USPP1EdWPmBQ7qYVi7NYjMRYWKnItX8r3f
IewOPWncajIH6iopV6DkOP4i/b70IB4oNWAswhJjM2gXf7SWByhLpxG4EZsamh3A1bikoYRY7A1q
1EUBIpdwjMxOJoPvm3e4qqoQHYrcxrbz3lzbz9tSITd50ifQoYLDPfBYzypfjcisk+PZfcn5NyHf
89XwAZ9i3mzS82/gighWqgPZorLYn17SFVYv55c1aE8xlh1nPO+6YBxcQRTpguZcGRjynqFztSAO
qPTzjl9d7CMdCR87Bzn/zDiIRIFe0zNqSb9x2uraDkq0s4k9cbZufIyI7X6sdkYlyXupRvQOuEDQ
9qlWrpokWSw7C051Wf6YitUDG5eOFPcVGAEhwukPV69zGXSaJJYZsxM7/Z25yQlMbB4V1cEnZktB
AzlaVxifjoDonz2IUvrt7/4+ondhb9jvg4cfmF8SO6l/86co76zTVDyfhxRucvjoEMEleI89ka77
DWaCGWDqZq0B2j6uhNM51PXqaUtMWabCOQqTgXINh1bi4VaYT+HP6P1uV0R7szTBFuRP0RT1vzfn
em0DAvRWDzwLQEt3N6f7WSg8kFSQXk2cA4r9jnlHESJUwzWEvkEGADFc/gp+YssVv9I+QKkUztIq
xGYhc5g0+hKNMEuNxE2ceS4N1ZA0AXupXZqIHpQd6PSzPPssWencJ8CealoOxQrnUeUIIq+2z59/
kPvsWIyi8XPKs6NimFyKukEktealDBoX4un77Pgm+Y0YrkeYrmS/Kfxtty0GvMiAUc2Yfx/GLOb0
/qV/uWucbi+UkzIR7OREk8ephTWHb+s6WqV6tLYjz7ziKpJ0yO9UeorqNupY8zl+wJfRQjf1hSLA
wWYc05RvxPNT5CHbZTVPCZU6NDx5LveVtDP+Rqi00T+07gyGOc5GsZeD4GLxR0CWnn3WgPkj6TTD
6PLnjYXXDSZhW0jSa8Q/EtZu4Ua6Jq7zSZIg05DzNpywssCiQzqTWKoCulM+pKwBmFm6Pq2bZ0nd
0cGGZA//ciQoijsTx2cZE3ur/0vTz9hZGwispiIOx7LsguhBRdX7sIiTfkpYxa0is7kpSG18CwHY
666PMEXHgBIgxC+t0ERR0B7JluimUowJbIiTYL6qfyNSzVBkU+VbL+AhPzIQ9FxSRRvk/wcRvW4D
pFXRmp2BQ2716r7F8aj6Lz+KhpXscK7aR1C9HSjuT7Hy2XflgjouTr0bUaUzr5hI9/n7dFAIa5hp
psqxeY7gI/20TRJFRNVvffVkBmcAwG4nd2L8iqRqtKsjU9rz1BS6QL/hLZGGfgYPBYjpXmTR0v3e
L384TPMFImIDNe6nBKmE9FXVKK0QYd/8NnUjn2JueyMZ4cM4zXxVAPAPZcNELqBbA0OwHuReGX5W
PKEdkq9DBb1FlCV/UZ/Yh6Ppwfc22aI4HM1aYslxBWR4r/CgHFMWBtfXfn+GPEuOptDkalnuEB2L
dPik+WppauCMCI2vk0E291jhHUQ3osM+g+yhcnDvgZEFmJ+NqIFHPRoEJ8NzmQoJpVrVX6bCr7DC
zkxccSOybV+nfXY8zbE4c56n/vjUq0NM1py2kULGTWVeGEUPwRlDR8NQEm5Z6YaQBszmHpiUxIrs
VB1VGJBrmrtwTi/QC0JBi06Q0+YFbqJ0SiRLmrxFdP7OJr1Ghg+XgcPIA4uigSWxNtggfN8De2qk
VnNkXF39zBAzbrS9mADhDE3QUMyIXQKxpqcYS3NAHG2urz2193MSy5Asfe54s6Deg4be5ZhJptim
gF7O1dRO4FbHu6MJETZrIkrRk5Sx9PdvWq4qnrzaXBhs19DjHRmB57tvpfTHWOFpAnu56G88lFFa
EUC9GMpmGBBs2FlETg64gruEVsAHg5Ny7t69trdqMVs1j/5LZhf74shPY4Muzlt0KYoJ4CFCRIbW
HfEBZOtuP0RRhIBkGCNcv1Fo3vOGVhflX93dVYqCDrTsMuefJhXTlzeK5PWdSJ6XJsa04W/2kDzQ
uSTw68YaJAavtnlPijcVH9e6uFT9399YxHOaCf0FVNpKTkyjCBpO4YYjKBopva2oCXFOmVw/w6qD
RFkZ/U9jbBHnfKcrUzTU6gLdSYwlwCvbRIuiCW+0wmPlDuVy3uSQCJaLVJ/9mvHSbE3ISOqcgT9l
5H+g0txrlaaOrTErt7ncE/Y0VRnxNmCCaF3KbMF9y9ljDvphfcdFNLY0XWJ+7kBcqbLSUNMlAnEq
tlQSfswHhPgI8QG1IVw5gTSRuD6KHt1EVC1GV/Ngn9WUbyy+g5HSIx1hngVfDiW309Txj5kM9ajG
Lhxq1CiI7qCZzBpskXUTgaIqZJmb9K3XWGy15bMjve+irAFm5lhtYEG40QwJVYaj1j2BDJHUEqB2
CyIXjjZ1RwlvVxiRRW3QQG/zHTmtHtBENVLLN8i9XYf6ZiiXFDu/1j6OZL1noMSfwn6bGCLu2s/F
t8j+Ltn+1r8jkpMOo1Gd0IZyYcMVV1t/2gGjpCC1YYV3eNTyOmbvLwJZ7RNXHD6VK2O5BEUB2451
F3PRkkvyo+V44qQ23aU2/LwZRgTHu0PDhPURAjIY5fvkSZbkRAX5BNOyQeeZt1XH6mEOoAR9jDBU
9S9pG/H05Ict9iJKuCgDGtLoi5RS+TEcrR6pEDqWWxTsgXI1jMhwGsi2rLD3uKSR0mrHh6lEh1Oy
Tp+5/ffsNMRo/uFDpzTTp1YzkW3J8LZNZ+o1F8cC/X5ZhgC0Y3uDEOo6ubWmmnu2qMUHr6MwBUJY
Rc201A2joLxMu9nkIABYufOzzs6d9B//Z3xD0vawdqhUXZb/vFbqgvc868ZFCAv+X/4JKVsvz0pI
7a8tAaFVMrgVrPfSyQ7x2h2+oJ1DZxtZcOaJfT8GSVgAS7jkqTUL9IayaXu8Ty8Qlw8N8kgrzF86
tcWK62hIURHdZLd3LIW0guiWdyMR29Mxbc/lr4nRWYT+21TnY8BP2WILeFm8n2cetr4Dz6yCgjjc
lMhTDYK8GsBnEJeVENQeYoPH51ksOvMYxGIFv2Ul55Jkw8sxptsdV6m7RrJ5UmBVYVAaT7QcmeXc
iZ7rjM+lCXFbQVFZYX9/I7vd90IK5QpXU7MSxOP+DujSCQeq93CP23RkOFWdW1rKFamLtLi8ZT5b
c++XxOELJ7ecT97pOhYSKiXvKl6fMN8uN4fcqoJE3N/WvIzJbgFuN8ru9W8zigJqivi10Af4L23b
tFSL24vzSWPiVMSK5jvatG72ej7QHPVezhKrUdcD9UbVY/i1rafz2338REd4+cWTNDcjnowT2IiB
VieZjTvdqcgV0VLNcJYa4h0pM+tuYUAHi66UzhpNnTrwgpoR+c8PbkLqrT3TvaRSIEbVc1NEF00c
RECIn4ynVw7lRJQ86F33kklE0pTW5k/VheXcEXGuJYHFK5OT3JNi+KMc7Bsl9kUMjC2AhEKWRW/u
VccorOtq2DIBI4Qy/401YRXXX97fVEOMaQxU5cZstTmKurdc/QqBvAJNhvm4/VMh+OSsMR6tJtVN
pqGgGnghCBxkwRli/zCdiWGwKUrBc1lINmc9prvtcHJQ30lMN6Rd8A9eBE8Yodn8rr4x1Sza3UTk
/qoUbzcVLUUed68KaHK0+XCJ25zJ8IzWiEBDcaJUfvqJwAct3XrYq5BcIWrDrg88fY9jD8hWhRPO
Vbxn40F5pokc29JwhnZCv1LvFWiwRBcWtiu2h9MXFHjcbostc1HR6DlK1EE3f2I0xqbvuaSX6Rmg
oJfBAeNxTl0GsM9UBEbmQUGfBJcisDKXkYninXeuT08vXdUDvmlYzz/MF4gRtitKcU+yFueweArl
e14eAqd9ArcBpOdIIkZdLPkiOpXZASsFv8XQ9ha09oxwhP1G6W6pmAq+w+vrkhwejK5DOlNKqGhZ
EQLJ4N8JoURM5BSQKoQB3KH8CGT19wI17JnXN82kWOKsBDF1rlXC6lp2E1N5hRmr+4WAZbV53Eob
MPPY67e7YX6yYYE1ShGhMponCv9E6+fuGl6J5eLIUFRdpCIOS1001sjBMKs8oN4nWs3j63I7gjVv
eLFOkEus4xUglKW9qM2Pik/9dWXIAfHarbSQNgzVeXQRWbu1J//B2s4iVno7lfloJiOZkzXUMZJH
FhG70v3NU6Qjk+RnJWShlGGvfPTem4BOqq/Rph9L8IqYj5roWrVMGXzf9vdrkvPQrN+6KbhNJy3y
pQgQGJYhMqmyuyau97lzmsyofnBmKSyqe/Xz09PL3E0Sy8b+knr43qQADVovPz6ExDRdZkgkSjIn
wGaZPQC48hIy/pTrjObL7KrSYJvcwgH9/T7R88YN7NnUCGQ5cEvNPvbQIzTCE9RfrSszCJrRHaeT
N3qMgJG7XYEtAtd6CyHvxnu73R+mUm1HZRKt1bmdnZ2oepjAMBHWS48v3cMTJ2fM2cy/excY+k7/
357Oeva+yEOCC+z5qWdZclj0vhIVrXl+/mMF4G7NsV26gzJW5pam+1yQ7TEXuBER/UJx+WRFWey4
iGgyjP9CWootdtfJkfY91C/cT2P7bZvFdgv0YvFlOPVasx4s/x7NJJIbnf6n7tQpKwvBYnQST/ER
VQcXIxq0B1+dSLs5oOohL7EbUSAxPCjJN4MRpRPdVO+N8aj2Fdu1OHWyKGtj/BwAVUj+OfKN8FN+
5UW6ur8MsPdZxJC2HQoOaAhhAYzDRabbTSFC4G7ME0j5dzHb9qmtUcQGyMhmEdGTbW5DoQIdm9aj
rgXZpLAl0EqgIpAngfEc1quPTdxQdubzNj1v3J4A7gA4wz/AHBqKGjP4V91Uc+xYLuPz+ldda1BP
8BC2TMz9IfZ4MRpYY2T6swhKI8j5hr0XGLK9XbbCzKxTw9Z1ccoS0A/l3KnSW5zJG4f0dMS/oYS/
SEvSIuzOA82oFDm3ip3bb4yCWQmsxIrPjh6cDGNkKb7SUntO+OPDn1nMBzXTfeNTML/VY/8m0Tw2
+cwm5s+N5K7+APIYptkjIezTfIp/MLbq5nIdKo+xH1u+jZed5wTUkxC5sxM/RvqNUOVrUo6ST733
Tn77jZ24Mp91zWbHlBlQ1Xub8dPHYaOXV1OOSWR8W1FzyKbNrewh5mymAw1gSkluIu8AxVr/BXbc
yFVfoj4HoSRzqKkOqFr71wTu4Z/PDcVXfkKqC+dD3UvOsk63o89tZhm60XbfHDlGWmgpO/jcxzTU
D8evltaaFmwsYZLsqPexfExcrhlD2Q849KSJ5zB9RxfFWBS5c9sU2GgT4/ImXA5SJnq8J/Sjyd+6
So+erwgTj60InBvirarFcX9fxmcYM93zDX5SfUz6vjbQCmjmpBzWB1xuA2tDni0bY0ZqArlMJH8p
9hwnfny+AJWJZHGL42Og8xsNxy/zmkktvV2Ge7RWxbvFXsqt/vxL+7/MK/BXltV/npKMGD1V6Qpq
O+Nfk/2c/BGDEIkPKRNweh23UOHDi9glqdq8wU3u8q2XscP4SEWNzX7uOsbd8oXumW4r9stQMJcp
eyID9kT5lQP/hbIQOtP6Wbd83fPgVVShIunAhsoDtj8aAerqxoOXsnprBmwmdjDA7kGM+/oe9atj
hfSOAta0HOld7IY4uuqmhlVMlK79fw2OGry1eE5HRFv/q09pxrJ2VyBvIwNyLzRwXi3fOKrX33qH
mhQI255DIWdkKgjg0fy1IwpFQyhhKSCoNgS0WPDDprssoK6ewy8Ttskq2bY5de+2KwUpIJ/4c17M
6Z6Wk6tLFiT465SoiRIb/4cIkQNMyhjEFVq2oNIqiNLR6QlcZLTlzyhwtceezLRCa/IZ/jsM/QD1
PmeQIQe2WAlikmob34bF0tO64acb2OpUrfCA0Y6laXPSdnBgIsYu7UkuLzojkrw7CpHUnsYWzqcv
oyQIhmN7QumIg1EJ5z1pXGGOUM3aBfoiDxV+biCGE+4zNwfmxf88KC0MUPr7mucBCH6SSxR0OSEV
HLDG89kk8R1Sw7vXBB1G5cwel+UH2hvc3YjaWfyiu6+Mi8L/pqsh7igdWrEp7lxxmep9nxaFr2lT
tjSL6LvmJphBgXiEYFQZ0EQ4mI5cKOeQZMwE6t3hQB5ksMcWE019zoOss/6451inTn4Y5O2ahVT2
p1oUboHrT8olgEyxn21KQdhAzy3gNDRUiNXP/G0J+sEdbbce+U+SndGYMeoaM3V+em3AThdzvvjw
XysJdeV2Lz2OskvoweX8VXObrq0Lzx7YLvQ1GXYf2fFuMTOk5u13NekX43fGOoUWP1f6cAfmNsuc
SizSI0LQRKCzFIjkBBUjQQt9LwEpOU7TgmXRjqKo6FqZftxmoxk9SBw+ogY7ii/hlKzxXF0XKhqw
Ueu2jji9IweC6EomilyuStWAv6w/nkN//j1sOzAhc1I+ps9Ggo+yEd+hAAPmrCLnyxnqZuJQcXHf
rbPrFTrad3tL9gs7B+/XEg9tIeGouY+mHCimw9b4qCyFb5PoTzMAAEg5QaQBR6LTIgiSCHBNcEw+
gPA4cbgbSDF4liWc9u6l4Q5Wm1FpppGxnJY+w0H+vHWjjuFF037h3gNquZToTDcSksknBL/MfuBQ
/wnJrpcozzuHZw8Sl/d6jqYpAmT5qd3fdraC2FALkWUU6QQwDqWfMDNTTQLlwKYxuMYqm75Zp5DL
sx0uNySYdtHL2U9U1dndWseYBrNb1m7gvz1TGeL1YBxS0sx24djJfs31XgoZK8BOGtFfz9tl5cMv
BtlGTMCHEV63cKKhkCO8KaRJKZoG5VgvoywY/pcLmLszRc6r6QdNqzqlpr95/a7nptGMW37bGBrQ
B+QdcRRa9jeKp0KRdmiKsUQRzfzlFvGpDBnni6bUMY7op3NckqkYIWuDPTBWkaX+fIIxqzYRTTfg
HuSVYkOoVNYnZQu5FyBAF92Gf4ITGcoZg+hIxKpJ6K9lBHK1gz+zfQG3qrEaoKI2C0b77gSJqKJm
tSLq/ABF2BmXRccyfiw1ngPU3oqTYUo8+K1sQH2HHJbCseMI/i9dePJk0bZvaKznCJt2Bkpzi/bS
TuywLI++5K8G6EEi2yQCqhEhTcG0ZstpheqiNg7u3+cciKiqOoBuZTbraJnfrySbIl3Pvo/OoMe8
JSzZQeutOeReUnnnVwakxYTaAlq0SkJIJsNGlR28vF8gjJTmFRayPaU2QMtJtxUt77x4sj0urTxX
KOxPk+hUZ+qIER2wk5qPNmXvcr/P87IQckEiX3HsHUeAtUgiw/h7F2GWvJNzBr+CdhP2L2rPq8Af
SaYigyDVgqCjVkXXslY6eIuCuPqArR6ru4uCpS0Ty/baOCeYky69czbYzx1QlvhcSaaF9K27L9Z9
fiba+PuSJXCdy7uU/5zsVoW8SsJzlVa5m6/puV78pXGyfc81+l6Yhb/bgSaN7x1189j3gmMfgVq4
wHO2N4VftPIgvSUwAJ6Ci6H4ns0WsQWJNvjt0Y1KFbsOVnRAyY59sLgnJ3XVBJKDComgbUpDxbPO
Q5/RwCYCWTGgaYXB1W6FCGC6WQHH4Fi8uuG3arsbLVeel3/ZRml1F2dI7EUcTgogSs9RvVRthx+i
33YYBJs9IJPKvK1HGWG7xzi0jRyLB5q1kgBAMNh9i97B5/caHbGM9oKjIAAYEBXp8odUuS6RVcnJ
MYU20/mb3A9fpc+em2peheF624JVmyHHeX/TdvEwmHzYx/LZK0ENhD11SAxHOm2Rlk54roslhUR5
qwcxJq6eTDMRbutH8v/m3dmh+QzQAK8yI6RPYOy6CXHr89ZItuV9qXS9Evj5nAViuWQ/KjvPNPu7
x6nX7kP3x6cC09Q2BE2SgC3rDme/3vg3FNeBonmDsCk8oWzYc8F8RaU7CNDRbMZsTEZQepGbqFO6
Se1nlETrehauXuwbxC2wK374pNDqbost+2FwmbMS6vxrHPvmkmZ5NPUMwnSDHJ2QiK5h+Fa6mlcD
nKmFySL1kTd83FD9+Gi5cIM/09Eqtj1X+WtGnGM3tsSDwScbJqTAHFD4eFH+o0/8yfsqVB4GhTdS
RZpbn/EltDgk8wUgwxnbiRslBsbqj1VJVVoA7Y8n0drwCSWxSuAu6QscFA6NgRpC023Sl2hBy6Ev
lKUA8941hvQ0y8fsq/9VJde4xBre5u5y15m7Th6e7g8kWlIUPzcFSrcvXrYFymuztK2TQwkyD2eF
1e4nKtUFibaXYughTuXdos8GoK4GqK63Q4LFM7QyZTAc6Oy1F3xsgWhUS9x1+a/NWDDcvjd2ZWi2
IA0UcMAGsaLElFHuVxQrYFtyN/QW5yXdArzQQpaNq8IcIfziFZqBUNoiptK1UmyM1RtPVn5NUpmC
5dFYZ9nHwH985Q4TClK/stY2MQqvX2dIa/DuR5oHeObSjnb9sqmgoqoNIyVsEmDjvg8mUluf9kNu
YnGgwy1pnnoPDs5ly74WN1es7WK5olJg2kM2v6Hv3FDK2v06P4IurqiEcEw4mdfgzeCcIVGmbO6+
bLTPaqkqau/PLhlKHv60IaNhpnWkaSbQ+CaJM6A79+BfplGyuybYHgJZw+SZRsP4StoRK6JjbLut
hBmbbaNDgEiFVwpdbVVz0OzT0YYIWm4bm+aY3W/T28t4z1l8qyjwJPhD6ym8IcqcQ08L2idwwpN8
zmgDI4fqY1Uk/eb+Ay1WTIi8ki+PcUX1j5GyKtniDGJEGTn2Mk4HOIkbyaa5BhlYHND7k1STzZ37
9ZQHVmw11jYiTbo8NiWWi3iq2ovNN3UT+mbJKFY/U4X+6ikPORNTh79cUqekxp1Xdd7d90Qttf+b
y8ODT0brVTfiFA/zI5v6n8qcFP1GcBJuV7O9CyIH1LmHEmB1SqSGR/uH9tdbOG692yi2aLKxU2he
jOKV9m3mZ+mCnmfW/VFFcpQgS9B88n57ZWzRJqUAHHNHtcKfH8CZStaqC7N0NasZDh+03Xgt+Irk
H+h6E1LJP0btsWe1B7s+kE+P771hSpAAh4JJShGEJ5mWEeEznvtGCSaJLMWj7QZQGfpMqpKVHk14
bQgyxaKG5RUoytOZ/mgr/Hy3xAMfKy4aeuxb/pNworY1jCMviiySrPDRcSMt/OlXVpsnen67DcwO
q/mN9Fzf/Hana6NpRByJauufTQ8oZtspICFNnQq1crAFyMtMY4S612BvLToiNOKVeskXmGHYfpK+
xPpyeCjtrmScM+wTZPzqMFJlcz7r9UxaPyiLUR4H0UHLOLwCw3TOaG8ZOcF/RFk7p8Oomk0t9Xb6
4CoXiFrp5fiRB9GCI8Vfe2KFSdx/qtuvV8NyRnNG6QXRpdGiHCmCIZ0BtVr+THs5Z3uA7012Cbgg
aAvwqmc6IhWvzRCe8jhcsf4x0y0PjYTTtMD2IU5WgDWdbaGSYmjE5PDn9Yh5+9nvY4PGzFH/W6Zd
q8adDzBoXylb2JgY8hETvS30JKj1hBqPAbaQVTqS3spL6dzVMc/9vJbjP4wtcxZp0FWNrC6zscmr
iFiUR/SHQ69x+IZLm9u+H9v2WrE+85uCylhL0z7PB+QXRwefEfazDCRYRznrR0ywZA7363GYaSIf
gS6wVER7B8S8jdEckh7KhksrSHjZHt5swrRBD+QT6/OfY4l7jmdGT96OBLl7LzsrULG0gRnc1BGM
CAO8iYb1vV3RMfCZK/wpNHgw/o+LSHaUblKcVxYqtz0azU68LZ5MA4xn5kOCwAv7vsRcLh84oJIq
US6XufUfKGMTAljq/qUsQOPzB67yyj1U/7qqUjHUmNttXO7ZUWQY2WDCRX7Nw7TG1+YalTRzp55f
FQXSkUMdlhKRYVWmuAS3laz91p1NDeVu9HP6FEpMfqMYzWJf3Rfh8pdMWRLcn/+zrl/zE9AY3UdS
HJ4B4mVAMu7d8FRKSaAJvSZDn7mXCOyEcbWUcXs35C+vPQ13WWZ0IrgHXgeimgxLkddy/Pg//xxc
sFI6wd/ylpw76FICJhZPB+tBH5z/erJCEMZ3dD80OiNamt4MN6ZolQjUiPYZjKmzyVnZeZt+LhQL
Xeg92mhDcki+ifQw0UxmZEszyDJ+LGqSYaZJu8NYnXaWPu6uUWd4b5rpkydsAPOItGF91P520ZC3
MJdnC+soujbqJdd8cFGbLE0FYD6eCAbjSTyN3RUxZJz/vmH6xGeszYfTjtSY2jxf13YJaHW0M2Ms
145VAMVVMsWq2nqqbcJLH50k+MuLHqxYEr6uZ2fTXw/oibPzBOLVF1+Mj5kcRkRJJVU+Czd5q9gu
4fGoojhccaT9tSek9J/+Cem+BtTWSqi8BSpML6O2tWkz6y70w0i96BzLJTI2d6CfRmcox130cDYD
u4CzEgyj8975hCWYt2wjCFRT/rCB+EyjOpanCCVeAMtTuYFBvsifSuJ1oiZZIc4wdp//kAhkzN7e
AMb8ngs6S77yDsOhbqxhOap4wbfieVSOnYHmJPqcxS4FGr3uRsVNUZsucS4AemuqDoL0nlMXypD9
Ckx+9nJd2DWFzQZEzBGsZKbmldJZxRGdcP7t8XvPT6UHmUqf0xI8X+aPSxWl/4jmlDJB1ay5TAwv
7Ntjd7/GO8FuA92IxKMSD2c0Gi58tjd4zdrTI722FPmN4HDgEU0iuArUon48L6cpsKg8usQNZ64/
h/qG9EuG58EhJHwK0Uca9+Pr31Z23hp63R/wYCZdjyV/w8daEpa+XZqHpqSj2xGxVl0WWlGbPO65
B8zdqfBNxsJfjtRov97HQ5ns70EPaH9ETdidtrMaBZhULDamcFGm+OThg3/Uet3VNgpVADjHdh0a
DYBma5hBtpJb7RRSOVhx7lSxENORn9RdCDH+YSrgg+/1rQ2VoDNwZ58OpffoW+Iow2cHgPVbGTvZ
8UNybG7P4bHYJAM41FlNIXQ4lSFf9IEmgaDaPoAHooC/wtZpxZgt5DNtuYFMfuuKFoVk+2QxAjjZ
gI59LO0PCp3Yx4onzv3KVHP3qAlub+BVWnpt6srr/Ye9fiQ4AWaKMyENA2VrYMH/ZukSx5hvrcpG
72gG3eXW1UDAl7DGpl77wfwMhlaAUiLnJyhgUU/U7S8mGIuM/lMyOu6CZ22GCglRQ95gytFAzWR/
16riXtV2PZadl2cgwi9ii3kqdhmE1LHaGS+e7gjHa4Hzo78EiE0a1iK6NTZsf4yAepjE4T0dZK84
dp1P+dDvh5qIDxM0MB7B9k5dyye7N7Is0h+KckXrgTZj4keCf5ZM87I6vXmrkrotjB7XzwGtDpAv
SU1z/hfEDayM0kSQSXMnc26t9r3XYzapqo7kW9PNvge+rK6z70eJX+j75JCc+/GmqbqiJQrYG0Mo
t9wdjOzbRj/uHs/8X8Hnk4BwXKjhRQPH8fR6eUSQFO0oWw2sMNPnXPoy+UD6xFvyTq0UgMv9OPQV
54gMCU81LsRqjEXQdVEwDiPQg8BNcr6UOWwt6nPq6UyngIhbSj6D+zSK+RdWU5GXHbydZebkp3Yx
GQqk1Rl+DalGb9ontKyp5qKdazWw2esZuLH+bZWUw/zLeN2Z0xXPtCWP8M4y+BkxP4u67bB3I5FR
ph6K6YVuAbIC1uE/IEfwTUM68rrrgO8XViRgKCFk6Pvy/gl9bo/xkl78/33PuGKMdO5eItizEGOJ
PwjX0w1z+pi+ZDdpFF5V+ZkSrfg8JTMzmPHlmkr8wcltjH+u28UFpEsV2mD6kBHCVKQGkKHfuVBX
OgnDHYDcN1fKaEIQoJSf+jRObbFJMi8vsO/ZtcU02PfJpRNEf2ZB7eOsuHndtPP5CIHAoFUAYu2K
k0afmEViMrIyYphOfBRbtVFNw2sVpXvaEaqVKgp3VYszJKonnp6UFgyhQ2oSEF0Jh9rt7Oj/V8tz
O0rwVfxBr6vK+U4G/6U53woKFqK4TeSQmXz+YKStfp8pc4Knl+mpXsyfiuZ8pwU7PauIY4RlEU+T
oY+/QyKqBqYR4b0SyOUD7abRTgOPMHjsATiRlONb4tCcQcYCpK0SJ7XQz7xk2bl6rJKhWvhh2RJW
vWqenJTIl8UAyI/A3DkgjjrVIchYwtKkLw2udOdNHXy5KDqEvTfbAnf/PK2KcFACPL4GvvvsGO/O
4PKrtenVsPf5MJYyMg1viuKJu7iYwq+Sw0kbvoSAd6zt/L+SLG+ekark3eXF6UbyOhG4gcgkr8uf
q+G0RtMI4HTICeAtm4zcNfGTH7xhuAqg/L8LXdrvfGkLCwETPJzfdreLa1FeukqvG649x470QP6m
3qwcv57luMV8lxsfb0RhjloXf7SupjhFEwcWQYvYYnsXsGEk7ouihvjTA9U3lNPGdHFXjofWVYVq
kxNLevRoZ4ChzwGxgS6YQCbME8b+5x0ekyI28RubLaMzCNJPIpDbSsnlqW5wXcZPaMVizyyecAiq
vba7jAH2/5Q65KsAQg7qsVYq3XmhlUg4etOm8GjZsRF+qp4mGIjW/G2h0n7aSZlWIVRzdgpdSVBx
kUNhQoRjJ78VexBN5Uz6QgASAkqzU1dIflf8i+D9ZgrKCn0UAGsTTx9nHt2zAAPgNPjdm4SBy4ef
CFHxIOVOz+VVg8a+jPB714by9G1bFy0dX2Cai9ysulgDRkqkTqQukeJYUdfmEflT1Q8U1nR/DYRC
gAu/NZpW5W4z0TTMC40vN75H2LKkyP+t63ilAcvE3bJVfOHgXYzBSfotNWHP//KXduThGQLIbR/s
LqXoMaqWzh8IhqN+ight+BD5GTHiQmxPDR8loUyXdoa6F5fhr/E1D94FpJZ8wZPIcp5e8VRYeIBm
GNDm4JI72cwfpc6qC7Rfn0EGZjM7DVPz+497LyICohL69M6lPPjga0ptiFNFMBy14N9qwAc/uuUq
kfoN4MdTxXwuWDPdnsHV8ZofyxJrgibyfClOszV8spAmv7dbMLd8ei3ewyxbScj8ZQimMFK1/kl4
5UBVG0Gckn03m7rlelsnoBNymvxH/ZRksAJUlNZEsA4iTECwWJ8UkuTfn7vjeznNEJvwEjlOnbFZ
TpN3PhEXcyxyGhXDCAYWhY2vTrM/6aJVIPqbZRhYse5wnhccRR7evfkY5q6Tff67wdHgdttHggID
fR+p+MQKbmttP11opat1JuHUzZTbEeD9h0sIeIIWWVUn1ZK+9UniSd1PucFEfh67oSBISwXqc6Lj
Mqpr95QX1vUChNIeuxhxVPUPK/F8VZBDloC+va9cCoq2EeVV8vLEuX/7seG+nRHfRx86MYk5TenS
19djj+MyLLg0o5CU5IkdMotcnxbC18t+Xb/C9VanwC4YsGbd5/hKQgIKJsxLsomEA+phT6fbFAUq
vt8EjDCFMXBIuaWztohaD1Pv7gsP9H4BIxpSrPoRYGEiJ0M9AGn7PWIYIw6+WajexqY+1Q1JyoYh
2g5ctyuBNPXacpATXRpnLC4tC/rZXEZ2+ha8LXJdX507F72JCHCIAECW4gEIkFSNtyrkcQGZllF1
zr5uqsEAJTcBzynLR5ri20tbCvbf1Q/Y7lYlH+ny4bU72qvFE48Kcmpf36p4M6+degPbd7FdU5pL
/9ivV+jjcsuBV/ouS+NLJBzIkD+mhmLAb4Nd6DRi0jk766l0WPn0iLAE+DuVci59bTfg2svAypC8
HOUdffGOHYWSuLP/cPZy9qTtXVF+ybYizzZNm3BxpZ2/DJ61qg+fqppO4uTWXx51NJWd+T/5XDoW
19t9rs+RjI1wzA1F1zm9O4fq3NMe/ookqsrV32UOC42hqZViu8cr046KU8wF/PMOAdQ9naGaM5wy
z8FCwtZhfsYfTNMDtDKsiMvtBEVwmvYU0L9TR4ZRf+BnoWYOPONmaizB2PmKIOpExtFKxKmXlivK
AcrtfQbMqgJJYJVN7G+XxMbX7JC6vbYksWDyGzryh5gDsVIm1n96dC+zQy+JnaihTFahL6cgYyWk
9PgwVA7/fgByYp/KXfllO6k37XV3Hrcz1S8+BiuLwPEwAT7CGVMjc5yIbY1pUs0QEsuSVQUXEJtI
+QQkDvKVdY46bcDXwPWBLbKZtW/x3TwsaVgdMIqk8//xmFSnf2vSw2KL5imJFN/MFjFP7XMvjVAf
/n+dpCfB2qGx4J9+4qfyNkyESdy8uDRTd9vmpx06Qrc3EGRaamHbh/JHcFELvj8xSNL5xva4WYUs
eaIuQ5cGxAOKAzSH8fZxB8YGGXkU+aECdl+baJFyGggZMxCLI8s5vyvlIPVYiivkNhqGKDfOPTiQ
8deF2zJU/1J15+mvCGPus3mbEcmHcq+Qew1j9e9QeePmk/kKPl1/AdAS6AbzFYjHG+oH9x0frgE7
YAAE/3P4/3p4h3baUUi+sKm74eOx+/SEkLogwjPY1uTHTGlA/h5QmlVS4YO8DM6IN+cUunNVe+mZ
8UXlUtcLBEzP7SE3SweYCFBiXkOZfYw8Rp5WVT3Tr524fi7+G9ljmUg+UhE6OrR5O5d5UPROFDiQ
JHcJW/bNxcjKfjwf5e5u3Ow0yMys8KI9eOQ67pTHcie7/dgLlACt4OhjnW0QdrUnJ39sF2bbMyxu
3kjN+FPeM3OWLkhb/odwb+eHorCQfpxQ4rPFIYMkpSj3wiYMYalaQo70VWXbtrgtGYfxPi3hhBdv
SfBkB6UwqewYVaNraqeylbTEdr2HztxL5TPcyIoG/0SwNafCiyaa16dPFROiPEskcyxUljZ8X8d9
uetevctefa4A4oCkhBWcF1mVlHKn10lp5dmY7v5hKnBNuVM0vbvnCrm0p1rkljTkXY1UKjKH3sz1
1AQkPXNKWUSDFslEU18Ui3+eUwYcly6BB618yStxCY6+dK0eRYOV1h667hyONlYGVCZi6bSFFojI
SWfhuDvyH/NaRzl4uVz1urJXAO7NFwDS+k20TRO3dVG31rjJRYf2MidlizPnEoNI4L5217p8TsGh
+cEugue3jQYDHxcfk/sDZkAcGpASWqlGtW83lsPN2L8JM9YDyxmOcD5eqxqPc0vkVvqW12ILO2eR
she2TrE2cTQhijzOnYu9viK2YXPTaNeJTPKkKHgk7KZM/WZHE1pAgc2ex9WzDuE/jDhBK5XzceHq
NtfsKaiYjVMEzI/2dNp3rYAp1P0KCdds09krGlI2tBQFX7qhdEM1v/pcJpXU82fG3YSxMoObsVkG
sJGRnlCpoFxG2DO2fnsr56K0EOsIg7RfBOTAWvPwUis9/T8O5ud3sEGeYOQfJ82012uAqjxy5/8L
8fouUvZgKu1aZOm35v/2rNM8JRrQS64xG9THNNTMIq72lapa4UGIHAPiWHhg/v7J2LPfyiKr47jI
VJ+4cY859E9TMnLpoYRkruuQUsCQbWd4lJzkx/XNRvcRpCfpG5iNXcqNKXBHdbqwVvBF38UZR6HL
DlS8yck8Wv681C7PNrKy/COQORH6MhbTX8YGBTUbah/bPFWd4pGj0OZ/WOGweXimpiWkpjGCJDvG
U9UKn5g5R9ahz1ovf9yPNhIYrNPotdJSnouXTWlw5wWPEcUN4v81tF7paa/pboeQ23amS0Ble8L1
wQ/9b1MTc8BPV08Keg17i53j2J3UVGdIAU1Q7r3Sb6ZBWoUSGA/wZ/b1ez30/oFpNS6zdzbmcfnH
we7kvo91Fe4JEjymwjonZrvDcOQtXccgITr1YvTXUUuBeNttJOibRsto7lSPHnBkLZYlZ/OhhUBQ
uncskKt+zSpbF13ym5/esMvlS3LaKdD3Dhi0Nsq/qkVJqDXKhyBHzs/7XR2qlRGT8f37WsSRRO2X
4iRuz1NoGGmE4G+3vwh1WbbNRorgOpRVNdKnn2ceVwDmNWIYqYNcl78rAHQbadP4e1m79aNZvuT1
PR+Wt5eVTqFTKzTu//4EM+YJyagkDNVMzkuYIopb9019crXWOPg6TK9zjwrx7GxIUNAW66yqrtcs
VUAUh8dkOuSM5mveKF9Yu2t6gfYkZnFMQtx9DbonUhNQ7bDhpg08D2B7Pa60h6WSl9azloJM1Rhj
JtncYYZIJqGbg8qdLPrdM+GrTuuoLzm4dqAh2oNmv+7o49KIWcjbR8tSE9GeCrgnzIg/6my05e+O
/t3Gx7vWRdEqNbjZHNWVhvSkNk90+ESKBA7lnPa6BOV+Jfffq8hyRZ9cTl1mspniCPcZZLbR506n
sbWGHc2ij2FlEFCNCt2ALPgYEsyEJpTAUfWAm33xqx8mRfHhOLYAsO1QBuhWnTQd6PeZP4jNd9MS
EOyzy9End01vP2Wd4FYJPWsGTfjCuuiYkd1L1GvEIBW3ZGvnChWMTaiNkyKxVnrySJETopHKvzIk
DdHuUQvZeLOb7IjPbpzCvYE9s/hogleoc2I4fU5VqijcQMRV/qSM0l4TqPmSWoexoibpZsaa/c1p
+wNCxHIxIblH/O/nSeeBAzRoht4LiO4ZRnT6C+QbI+HjxEM4j7eNV5eVFFwaI074ajvl6ZvznqQX
Wf+FMMyF28HRVjXk3FMO7NMjmLEW2NAfNBanB55SDIi6jjQCtBp5VFFyxcwAp5zcNOCdHRc9S+EK
JWTkE3PPMqxcpj72tr62AOoDeQYH7GfX1jbgy20HCkC+t5oqAgXMhA+qADMR4gbc3/om6Phyo9SJ
NEXjy0+63/e1ul1DJmZUgiQRnQaWrE6nqU+8vQZVZEeTtHFj7Dh2oxyg8jiaxi3Rpjz4emirXSec
+BE+a8JhAkH2b3WwuRVKt8PQ3N6BRKMX/kOnNzxiSv6GLM5kLDXk0nmOOJLe/0EokeYSDDaWJiF6
ZMpNZFYL1AnJQtV0cUuwdBX8tJc0bVg8p87FayPJolTOPpcmB/dJWJXpKu4ib9gU1bdy0L+bMtbD
7Sww7+e/ScqrEULbleEWl4yn0Hk3bd97b0G2aarLSczypDwztNGW62+kled290X+vRmhqZDTU6+z
lehhuaur1LiF/nFVCs3VSZdklswusY2r5FUzAWBOGm1Kv+bDdyvHftZr2hk2zy7hHIbBopYHH9Ru
x9YDVxclo4qMqfPdpA1GEwM+XIdgAwpgzFH+DpGPHOGkXVsTdgdTLjjEkjCrfqEpbd42QqRL2KDT
kt2KJGCdenQj2W3or4wmTnT+oyEThQ4xcg6+Gga2tDKDPV8wewkbXAe9tyzZ0lPSeDbkhgoX04Mt
fKtMiCSdQAyJHEqPYohRp5NPWB1z63DzyGFprSivdPLp8jIkvymN3Q79WCmxR2Ikjs1HC4hCM3Sw
MqEvT7MPyD9TRnonJ04KiWGEDG16dJ71Lt2T6tcNf4HdGR95ymx+Edi40QzeXZWje8tZQVxpDc9X
2FDj8X42CZ4UJH1bAYERAN8xUH3koMhg1Dim9lHm3NZtY4HBsOGcdBZqSVo+cVSGNqOXFDHNNkGz
Z7IXwY7S5GYlZ95spBLgTVS+TiWvEaKTKNt6M9Iya9JA+B37BWU+wkzaZD1+2KKs94azNkZcmiJ2
YrTQ9M6f4AcNtkRQvm092dfkNTPbpj4lLCXxWKT/84V7iCl+4x/Hkkk3+PuDjc2tYeAQV3C8BWZC
sPBcpNSGSlChcKdGUhNjRJ/CBhYLY6S8xeNCcrwS54Y68GNw7cY6IwQWIZaYGQKanVb2y89+f0yM
3M/gSnHh9662J9Fo94dnp/HvOGi6kIlpf7qzg2Ajl7KAKmTTvOjFV8Bok33JSFCKS7R3px3hUdsO
CQoHhmmxPoJvalXo/eFGr8X7IiUB3LSpNwL/Qm8Z4l2tN7UAPQ94X91gXCWcEBVr44+IMM8I6OvX
EkK5EWGh/Hstjxg5e5upN9z+s98mdgtFWS9JSqbsrMWerZ4FYLm8g9+NqFv24+tLWymFguZ3ITIm
P4mVdUOZ2WEDZF/Ct7Fss4J32TrAzuXCvYCBx59/wXc/CxikjjKWZ/8j3ZwfnF8JFbOSNmgqYLAN
YOEgPtiWZcsqcETUI4faeB5errlNNn3RLDRThRyY9n+Nz8RIB3NrqHwoQyVxBKCEQCu4XovZN24g
VvpfPWYKEQw0NcCoAnR2w6t1+467dgs0nLAjB57OI37DTCELEaN5FWlhxrU/x74ggUzi5+k47P94
nrrWC786hNaT2EM7O7cCbZwvk+wVeWpiHXJf2FabAQKVrkvx6AzZ3bDM5BFkv2WG2KzS2EJlmmV1
Qc2aGCGAApXQrbA9dnHsE3ZlCFMrUejt3Z5QsDr6xxaBIxv9n6d0Axd1BK6sLuBjIt96DiyQpTJu
k663n6m/e8R3/Wq94/pykXUand3x1yx+p/2C+UgaiITBMVuC4ndLeQ8pJes/QJ88xwqKRpfXnvOl
5MOCrXs1NhxTb7Vcun75BB+tkYuIrvawYDXTKNLzMRMs/XHn1e6LtrMsFa5Y5xojshIk7HbBFMiZ
fqRqDBBvBNLgOdc3B97egazSpSqAzGEYmL6qjCgYIMIflnrW2lKkrBlDnfZIZzeCQeMquYunH1wb
iVev8L9JP4jl2ti5N5BykDsRZj7DPBMt4PehTOTlavuMbRaOcUg0ZrEEDR4FTdDR0fFKuDHMe8Gz
gTnyH7mVEuZoxhT3VREa7YHwmbDM0yHZ+Eey6Cor/ZDYCLUeoLpPuyOzv3cRXLinxkiyaMBQuiEO
dWrx8e9pe845VRilAVV3W+f37NsqjWL7dlMAlEEYqYLU6WdV+mcBfBZu6OPxhHRQ6x/vArjRKsOl
bane/5S6kzcaaZyp61Qgg9XP0G+xl+ylbhIOySaGHEErNKXzxpk0BDBKdgmaSto1eYNT2VeDGoYs
twpB6giCY/JKDbFQT00Nbrup21hGaH5nMXDYm6qKqHcbyEwPTU6znr0PeWTM+Nb45cAN6b0sENYI
aBrhu/kkuMdKEqZIa6xAHafLY/a2VUdoxl9L+r+uqYqvp8/spkniskw5xOChWk5wr5dPZ92Xk6tH
Vq6/SfshKaGQtOc0VT0zLu68604UaAVRNoxKxo/Nxb+aT3qzOdYHxqx213RlaDzXgE4KTKYRJGZ6
SLUIUkzCPig702Nue9YqLXB5Oymam9QuZt394uL4Sd/jL56KzCuKkJn6h8nzbZ+QtWG7crKjMt1g
tYwCmWobLHL9ZHTDAPX2HUqZsqdp6ohOpjrlBbMvVM/nJEjvO+zHvXgNz4Kh6ak6tzcyFSqkv1G5
eI0HTWSIddl2e9g28Hg3iNZi+CmDojuoQLbQmXyD0htgyMuKdwKmSbN9dG8dZGmY9dnzV/q3HNQs
sH03JH73PV6+VBIlNQ4FK4TxgSxg4QMBOAfUt1AaudWjhDAUGbXws/bPkYcgneTBWwa+MKuFaZCU
oVWbVEeVja3qCcg/hkk5pbGqvH3hWLTJ0xNbZB8IifUbkwSONgCJK3wOLvmZaf/pOKJdz0k3gkuO
je5ut9LLHrwQiOcUOy+puA523TmoqO/NP8472gIcSOcZ7EWTrNfLft9p1c4W5Cbdy4cO5eyjcLU0
NsY73yhXoygFxL/gLnoW4/eMg3rvgMDRo/HYGaQLwc7/Owo4/Pl1p+q9FG8IWiHIibp4+Ai5VfRH
KhcFkHGVZkQxJoE3NwqxViMfrOw6J0/vim6anDtgStS6wGW1fbmt3QWJ7S22X4ORWkx9tGVvEHr7
Hkv1lkCO5Tamk+5XgrGB6ORKHpVcYwG9oAYyQDVNyuz1OXyKYJvxh8CECwhrbefsnPHpuXfgWo5S
Jr7tvDj8L5alqRnZm4QOzFRyCfa0vCaDnn0vBteZZK0e+/aKCk1QHnz+JD7a6QLqecD5qiRtdVte
swM++ZabutJpSg3GF9nuAMwbqxzqO4eKey+tGHgSlmlq7Sq5ZO6q8du2cNws8TaITudNtMcnYAHz
EcKBGDPuU9P1Lq0Q2qmMOWzHP0Q4VMLwqi2wc3H3JB3nYtIph2jTkHVTBaek1Oa87bREsLNGKDOG
LoznYKqvGYxGvPdPuFlVPrHoKSEiGWQzeKpt2BkhamBXl99i897FEnYJBvpwrQUzmQ5TUMiKyss+
dpODBJbTeeto7d3Utkwofc08yMBVsIpK3e15Ay4ZnATLC0PxxGu1GtI0eKJnHDZU4Pd3Ea6T2Prr
3f4iKYy/G2Mj/vJgl2i5iXqAH2Tx4MBKEhUM9a81rD/XKMdE0xMTw3NZOxx0fbhUKleWqELvgAef
r6T7ZnmcxLHS4zsLDrVxL/0h+Avoxkj/lkiJXK49TrwYt77lg5mJALiemBsAxLcV3QVgbJKxTqwg
65lS2Xb1h+k6mhLscPsIC1g08BUntnQSPOMui2/7VmazeHIE2mqH2mzcmWEainJHIu2YVl2sS31v
G586ct92gFy3Nuudi4pWNJlqkqZqkEaIjQnDuFMoPAkwjvdjajrzdBzpHF93vIjdCspuRrFOlqHY
xkarq2nHH3n9vQgSSyjxUUwUDds/9VVWGoWxBEo3fREobRvj3Jr2OfgHi4XzFn+gyTk9HcT1wAJd
/J+xd+XIaY++0zdfPk+5JIqqfKSKfRm5jLjBRxsNVHcMm7lRk4bSBX2GQ893OIbXegkDmz8Vhzwj
aCj9Y7nYDA0jb+4Pan75XVHTnHiOBq2gTMqMeeGMla53lnHv7wr8klciCKcBA1X0veFNG0F5d2ya
p6OzzeXJTZGSNo5FnydYLimX/CdctfispO8CGRd0OCkDJue2JLNoJouPGx25IEUHidson82c/rMc
krZA7yts+zY25xKN2OaNDgu+O0tUianhPYF91rvikTaiElS3BMxsjzCDN1RuOVtffn/gkKQ0ZOmR
EqHenE4ooWMzas51nTKSxQK5spqoSVN9B19x0E5btFtNrGFNGhuBRtVXfS5C2WvwOz0bF9Nm0TAh
lC/PLLEd/uvspJrY3LY/cW2PVZjx7jViHLFx7K7pdru+ZFbDXs63eyCc11NLbtvuKubv+c/JyfGk
t7zHffX4i9KhvPm+3aaw7UgbH7tZz8ixFy80rpItQf1/mZhPw4bXQAkAi/EW6s6SO85a/UD5DDnd
VWGJj1pEpPqKD4F2ZlFU38LF8At/W85STahcnntABAA4ezDrjn3h7TYDxHa6P3NUVSE2tHdyrCXo
Hk6n2ijm8bcrn1wZSqRJextYj7T+FhCjfV6R17S4tU25iIS9/LaVtHbC4V2HPYVHg8yGxru8wZwp
aD0mLtpDuNyNueLILeBpVz8gnFyRcZ1qh8t9ECaEumi+nobKY2ocJOI6ug32u80PyllKY1SjMc2F
l7ktgevYTwUocJbmQ+twrynz2MV0wJWTRcwAftyiolLMU5kVZb+d/XXyRCXudz9NAMIBjQMYzYyp
LzimTauautH4+t09v5SOk7x0TwHyIaWEazHbXybV2zq4nzmn9weNyTtzvlo0tq8jM6aK4+TwG/+R
WqAZiwbULmxk9PNm2rD4+h/mtS7Q2USz/SL6vFjQ47KywOtTLDSyCAk3oBbh3g3P/TwWeXc0IiAj
w5r6zsHurbwQxb+6MxUtlNthUzRkUi4jZzFo2A92mT/plZndzWNJK1l/5/C8opb0biXR5vmaZqwZ
g7qpB+B/aVIIgCDfniBRKxhDudYXgfoVDI5XGTZtsS3YG1qqDJnsY0E/oEXFvSd3udjI+BU62Qax
qIlwzhulvMnl/4LEfESdWqeQ7STSDIQtR6xI727OtRb6a8fd75+7942Imt+PJ29ATm9Xay+PG369
1o3A3LZ+fqLBMdtLlZFll09YWNTBerzYJHlM6lDy9DOWjOWNA4Fp7U0IrFLOMAhOt4P3o8RrJUeU
0Ejuiql4l8sZTx1JppFZqoY6v2c+YliUlr61uJ+hZ4dL6FNT7F/uwbYM29NNWglKebVXRKSNeh1G
R8K1+b7TgvN+Bz2jSCCRt76UC7eEhoWEdI/3Lm0VX6Ero6vo9IhF3Jj1x6zizm9MK7ITzr9ssxe2
0/NqbioAoDquPEww1lfCwibwAqMjds+6ieTyyO+xxe4MScIlMYFO03I5EXmqYFc+dXj4eLQd0Dme
AiRBE8V1un+/cB/bO1MMW7JVQal4raCpZPD1RGEkDpWqSxMlFs7gLPCXb6k3aFCCnTeiTBTNHFhV
D2/zM9Qqzppy5g1hmv194KAi/OYiEoJKlTz6t/tQ0f7khCifSgx+DdABur+6drwwhvaeqo0f/bDd
DqQKncWAXL2ZWAY71sIltlkmhFTcd3CStW7mdACFmVkHlGst63zkTyJeLemuaoshS0PRkIQ37rXZ
mNh8I+yEN6J32gcz4bvZB7f1BwbSAUlBZFf6YvCArQnXq6teyu/k8OY6vQX35tyEs285ZTQeptKI
xjMIVHTc2cXWIeEqx/MHnt41apA44wJx36daC/4Ck1OgdUorhH13ltoz1A5e40eazVewv9myISgU
Q+Uzqc5tFXlJxCkmJ49KCjJx2laoH+pKXpNUQFC/GL2XAiH8fXRkeXX6sjz+9YC5Y9lSfUEyewp/
ndLJybDCQdaAsyM9PcfGbTO3bGyzl3VFNEU7pCBBk7lRrkBE2P+G71kand9Xu7Gd8YRxKmAf9gGf
V8Z4907OapNNfVKCErevDvizWodGobBWq2tSJrrqKAMQfqK1Gm1+cym3qSWGPrIqFLBnMZv5m89c
zN94qL1/zSUb0Klp5zOq4xwkPItayS62vjvfvGFFL9GKw8XIuWFJL5rJK5Xf/qsCQfWUxvNexJtg
/d/WgOmxFOgsO3wm4l+MgSe36pd2wHqkx8EW6CsOCjgk+3iKdE9p658R44QEg5gzxaCWPwGQwTKX
0reaWmly1xRIOFrbdqYBDft2JUWg5uESErX4OJeMk2CsErwuYr/JvHHdNxXRgbc+38/eDSfN4wZs
oWJxwznKiT0x5NtC1tXmOoPaiJzmyXAt4/gIuwRqLlmhHf+Z1DL8xBLlpbXjUNPRYIDSh3C3NML6
cHcVCjqZPQqq83ecLOrbjXxgKlLH+vDlQhKWZKNDR/FPtvDdrLTTd1aJZLF7c8+DZRg2umim2EXW
T5oYXdbann3XLj9P27tHYJYgCOctnrfKaPcd2PfAKGoMZIlOPVzohvIkNn4viZut9NHsJeSocY4a
4OFQcAfb/u6QLEYp+xR+MPNlLg3MIjsIZDpByBZEb4tUulKdazNrckZDrsoaPvAlgE8sVCeiZsVY
pFQieyTJ4wwjNDNkRRU8HY9AFE4qThyP2yTLwsVMnnh3KWm5sYyV61PJjrxIwGIcVvhPl30vaZzN
8ux1RAwJBi1x9jqG27A3QHbeY0pLmkp916ks1k8bG7MbV4AYinvUtnJ6HnwM6r/fhRmladzgLkRh
P4q+QE0/YLL+rGBqYsLcJtQhrqx3/NZBjG/lttAMay0f2scRIU3G945iGbT0XNbf6yZTMT2W7Wnm
C91aZPIR2m2iyKAw1xb0oeJ3a7+eMm8Oj4nFevXOLvL42er+T6By6AjjbUZfX5yvw3QPxSsX7Sjj
XHcrqitb3Br9aOVri9nAWAFeObpIkXOnnNx/YvTNuqK5hdVBozbtgaZJG1RVfaRo/26XwXWxvnR8
opir1yLlczcma5gyCy1qX+p+QR5BEA3w/4Ie8P788ppmnaYHApSriUEaKwYaLDbxvqyG0Ha+edpf
FzVyXmiCLjEEW2VRdgWnNbsaM1toCrWe15OwJg6aLOMFpPHSS1LJb4DfhoEft+y2CK5NckIFJYeu
CLUQsFR6KY9trHh46RgijivZv2eWe/JN3t+buAeiQ0xGE4VLc2SPQVavzxucOl9LFijzo9mMUHJ/
Ca2jNyWFxfIKzXYuvARNAj21JQvFqfbu3zgiGe6BaCiZKp0TN4cUJAaWUYGxFlr4lqajmPu2Q++n
36lZcIIvgUbbk/2D7sgkWfSfflnuYnaI4CTcK3C7V+TZDan4zXa2xD54w61lHVDEbsz0tX6pMzmk
RL9mrASlZxsfsld+zYO0ytywmT2hUrfKSK8vvYHj7PW91vJKt8aZGenGIxD4p+i9O3lwjGwSwFSy
yRXKUtCb2zXevVOjs1raxwNIxbLQzmsg6mSx3tPgeUPEGHdACAlv1+9z6H8zW6uEJeoEM0/3ltkg
geOOH7OLiu0YS1nip9PD765X7UUZ2THw3LiGCXY/BbM1COMpzLEVS7YMW/ZTHaUgofij24DlCzCK
VWb1Ow4BedBZACbBSHOHK9VqbPjpCrZxOYIKpmf2GwRZmmDXgBNq7bZe3Kaq0lQPV+iTLua7YNVm
nN9qok9RvcmON90Q9ygLft73dIR4sU21NMa62MZgeCPCcBWnMJmjkHZKyV+p6GAlbmB7kFdaS60N
zs+9JzEnYzNM6GUM+j3JtiQ26rRkn7RBxsyITbTHj8X5/MC7Si6NdAMVcFUnSjyCwfJD7HmjfiAO
/8V8JBHh09qW8CSnfisZ/mSPk3Bm0/Fby3SUJAOJCUwAe5Hm5GdTisqrpiXFt+rMbdka8pQ+QyAe
6A0yB+yUn9y3znFGRlTvSobKAGdmEsGHGDftdWH4u1ntKnKtfJRnYPnBix1vPVKq6hUAW/WWvraS
7GSsfjk+o7cugO9gAcMQXYHXhzrrx3XWDhbEfIuERekEpZFzpNQlHgmGfhM3UELNw8nBlaBu9E1T
i2XO/2mFE3e42lG3viGKjto7mr937a9TCmQKwR1yZklJMxzBZtWQDEPWD5n1HYfqzdyNxwQ5ws9/
GWC666v/ngSv/KidDTr8NOaIxH+u84efgXAXezfnmXw9yXeWzDhTU3zNDTZ3UAezx0JSkjTilWjV
tPA+Remq4wF+JuFoEn6hIMK8tLdltKo1BgLtlFpMZlr6Tt0AGZAsnPpXbdPpk08T5NxPKp/CR9+n
3Dq9xAmvInD3xNxcLmtpkBfPd6NUKbPwFCq7IK2OzLUPHn3/DfIfvr1r6fZkcO3nzMmVkM8axMaP
oU/p5FRYP5QUw09LFZdAPIyCO9bhNQTEHFuexIRBosrhDvOUk8kAUbPyZI7AaqH9sF6395/ZVtgp
GaYjyR5vPGAP/8dpuByySG1uTRLklKZz7WOGcWXULcgWjPizdppwYeflb/Ysg83lFnAjQfL1eNfF
sLUN1W80gdCeM2Hoa+rtNJbiEeuN8ROw2J8SQfKx52aIm1vonr4KGm2tWtGrrZSmEIN0isCRsCgE
n4R6U3E11YLEjOjYbu3GGOWHZc58b2xFjAiNEU6MFILsDeZMeasdWTCeZCJbaPjlr3CzzhqpmUhf
N4nlxC0JEWTbDhldEzfsNetD8CMl0yX52ra2miAYzGj2qApDRUYx283MbfcbGCL/qL96hH7j7cO/
mZfRqc5MCkFxMZYT7lyb73gsqDQIuA8qtLw+UGnhf9lIjoM3EASQKqbmY+6O8BMDpORaJeXa3WrF
+OpoWjIrLxyQtxfoE7SVHh5X2ePhQN6mntVZkecr4jnZ47smz9Vruw2J7s7VGl71BlovjTS1PT8H
MG0MJadLaa411Eb7WP9Js+BatdDs4fsQhk1UGAQyCp3VzHFFsYcWIXDzHIw49fuL7kl+qL0NLN+r
BbOvo+r37mVzcjybwL7yvqfjif8+WttqT7ICH7cX8QDhRsaKxI8b/HbbOI0xDAmD/AQ6EHqJ4N9X
hF6Y5XHm4QdKmh9kVxE24ZuRgAf5DT3PMZOJSSeap3FA8YJovqEosyW6tUWTurqGakbd/wPbKQIa
L7aXHRjQdfgQzCzc19u43bJC4wDYj/SHXQL+GfgXhsCzooUf05DHPJtpfNpbr9XcLQYi9UUoysUB
Nd0uqpyKPsKjGGm/cDrl3Dsv8TjBS4XMH0F824NgklOHOrAM0OdyCdi0Bxbhl+jW0vpB4Fp5Nb29
RbZZCaLthrBIIrkpqHKQoLYP2HnMDpe2AeEnAuBPyQkas6BzTb3F2UxiHGFc4hDLd9evZ22VCgI3
kRjlERY7sYPDBJ4JxPNHmB2X5HnLlc8H1Wzm7kHPyLq8VlfJouV/+X7xxwjs5uh/vrWMDO8GKPDn
K4T3JVGc1WM4o1r0wYvTipo5EJgfgTCcv1EFSehb+Oca2UodMYZWc4kdTDwUBCRM6zcrhQcXKwKX
TVNb+uZQCbnEn47hE5RFvjDQ1KWnTUXumxAR2GzghT+7N5+5DA/P7WfLBqJ9dLSOg5QeYHYR2Dzl
kUha/XEDjWOW9IWVhe+HMsiUl8OdBVvyZd1GFmIJNZiYu9qLj8ZFZJBGG9snGKpc2L14B3TIAgty
RIBtRTQJZDdF7OPL77r85cEs6GyCajseHtMt6fHIjQs0eSPGCvSGKK4iZGph52O1DjjkSpbyLc9C
CukKhIps9FhY9YsvxgwVurOeipMJQC/fHrI+PkSJLf4GCblELNMKfiXrtt4LlE2A0sdmy5Q05M5/
PgTEq2MoDsGjeJcgPcQkz7pU6cYQg8AujpFI1b0GIQ7RS9dCUbsBTywtgqP4LFZHKOA1TxiaV0Gs
zwYbM2OriWzYe/jvOkx1bJaCGoFCC7UofVYkDbc2O+XpFFMytsuYFsa4l1of3ebv50NnzE4VB4EF
S16tHQ6czKMuGujLq3Ayx3oIqPDofS7DhVanQac0QmfsxmwPW+TmSfOte96ReOIwS7a2LHyWLuQz
XQQu8OxbCdq70JMpJLRiTzk35gINHMoc/DMcYZjCCeyaCZ1PUWaUBAs8NMjNsUsNhZvZ9Kh/362J
5gE7x44hwW1l0Z4yrpKu7kxtkJ45jhRGjl5SueDOsygBur5ZwR/0OePBQDV6IgCzaTpCWP8Wiet5
vkU39j+5+VESeJl7ZN9BInLpAvH58GFB5Q2eOheM9BNzLZg9ZOIa74w9RkoiHyUizPBDyGlywY1o
zlmE6+IpwXQ66sC5o530m+GsX4Jcu6vOa45xZLJ3PlDLl8WenE0JBs9Lo9U4czigubXcJmFXlr+D
obnsek3jRI8yGT+DuYPhh/iFcVnjyf5fdfzzjgQDW6+gLKT0dhrAG/o2IC9F3kSS7NXJeduNkVmv
hETAIUucO5x4204yHE/uxJKjA/kbkdounRSFXtuwZs/5+V8KfDVlk1JWXORJakoC29jEPFMH9AVW
VB57WCJ/SKJ2gMD35ztdDBNPB+Rbk5Mhy+vHHO/PYP7THFCe11bK8F25X45Sqi2b3WeXCrAT9Dlk
XzX1yyNB1Tmq4Ieik94hDzggBiqE/DdvPele9xPbLYBWHCnnsavWGgA06aH4aiP0VXDgCCbcJ/0g
5XKzN1GUc3NW8ouUQ/Fqs6jPc2FbGKJSvGd0fWP9018dXw86RWBO48O1f7d5Jjmsb6pTVXGzEzuv
nFK6Ba7DC+Qiwux0xTQIUeUvvnaQ/pIDk4ExfQGtAUrgjzxeNTM98loxiUBSC2qhc26egfTuR9Sf
N5yT1YZLK17SFcFM2mkyUo198IMeVgdeS3F4RSr8cAX+w5ZlmfYUwvFfk1UATMMMtdY0c3a+P9TX
z0ZlqXp3DKQKTJPXAHzK8oJ0ahlIJGvp0/sUZYMqh25EaISCw7c3ULyTpiCBouN9eUkkYK5GN1ZX
/fU0xBMwA8jJjf8fcKTpPyx/3NcGhK295IcD23jmMY0voshDdsOSLmut2EnzhGeGCxCkzp4ZxzDN
LCAPKt7Xsv4yiGm9rOuX3k5mNWRNCFJmIPi6MPpOVAo5dAGmdkgnMrK5mpa2sMlvdRow646Bn8w+
qTNz4I6U5rnAp7kRxdYa4J4Rber/ohfK674d6yO60Qx41UXMLur7wbNFr+djPABieD48dnxFD0e3
b+WrSOaUU5rYvbUQGzOlb4m1n2RXFd50dgXlnf7LLwe2LkPYIPGQjSVFtLvS4htC4y5dGEqDQUBM
ZFP/QOVUDKXLDjtXZX4Dc7mDuROP4oHQgCxCCh0MiZ8298yDror6Dl3NMyTEahPPE64I6MTncZxF
+oj/Ma8TJ1BsNanUl2/R//oL9IY5NCKxPBBag+UFmxj5wzFVKaofhw7AwXjeF3aZjYWVZdnI1kC5
Z9YpV6fWWQVeUL3nUSdzLrxWZ+DZWqhrMp5ZTpmwwMcG9R2ly/EqhwldhPK+b6esE9E71nnXyF9t
fBW572HTgXp5/vZLQg4499NH/rVGK6w8vYlbiG7K7PrIkEgjrEqEaDZGrwtSK3YYyXJI/weZhd7t
BynINCH4d2p/vicpJ7GqD+EYeZV7JEiVoPZnzjRn2+u3mWOIlsxskWrEztNYv9B/TdB0RXITNhOx
UjvTd95FeRO4qsF4rBjVq9gxOoDT5Sx4CLmMEMmb2ER6RixfSBIMYJ+nLKrIb5p2Zszk5W3GX2v7
dQrWq3i8o9qLsRgUAPiGSzpfd9ZA5SaKPMaaoTppJ+OWKYZQe8sFLHr9UbSfpse13P0bgig2rggr
MxWvemqRrC/UG3FQ32TGpeLRlhzQopfBXTzENa9rYY+52EUkMSYLqGlu2DmyVlFr/UresaVcKQVO
2UlsWESfrBuVXRo4K+ASne6AYysOzN2CNP/VT5NYQzt5rimCNiuCx7AaaZAMtQImurP7EAYKU/Kd
kE3pAqL9NHvXC/f33fJNzmNgT/vSfBiv4V3eifECpbhCKRLUW5IDVdTsxMUwyOTvtpO+7Nmmbjdf
Y+teLnNeaMhNKEHFZi3SpFglfBJ2ljfQtxr2bdyC/LIOCMxX1nKzYn6ZVYj4sjD4yg5LJcECJNbY
X4x29hRajklP+uFZqJUQkWs2HB/aP16sVAP3/9AfComPBajWOp3Kta/rr5BhRuhW3NrfOckgSWYt
s/qkIiVHtkiUNOz2YQT6k5OhRIXKS8FJ6GwRplkmHT/yjqy8dZBJpFYc+dVjoyNAigVDuBemX5Q8
R/36lRT9mVkncej4R3NenZ3tNtZxS4m68Flo1BSOlHjUmij+TPgzgKv++giWx6amqyz6rfy/LE6n
OAhzYPGkERhbVzx0RAb+Y0D6ZqTIiqLyOpUnzrseh/XNbbhcTBsw+3lEz8mlB0nE+BgtLjmyMTYG
zWaqU5Ag78FOBB4o5J0hd0+pTCrRu0I1vttRlBVJmZySgNRWCDt1Uuqg7iAlm2Um4ZJrVDYmVEkl
UuZo1wf4phboLad55hm+yYol/VRAg8HkrMZezchsv7WOAfu2WshMnmnahXMEWiS/8QpjcwIo7/4h
95odAHQlKq2xSJStVvbyAxKHL4bVKRpVeIicFLci9rX7833798wAZ1GtZo9coFlTKW3TKDldheum
I9enpX1f+05Vw3nG6lM0doHsLNH2D/4BKfY2jp1R33IW4debCKPEKjS44VZlGIN2iKteMQz+3wth
9lnIghltb7LUeCr7s6YOy5Mb8OMrYA9lV933iyO/3wR1vsl37s0YJTEqqMCnVHT6oGmfgx1HyRgH
fy5ytS3g08YmbOwWZbAQqhKnGZHQHle1r9Giri5Z51ZS2W+Y9UXkuPiDFYePY6k2bmYS3RASylap
E694iIaIIhzv3hFOEXy1z1xVxDD6DpAug8R8WqAOlRod+R7eq8p1FDH2m8EsYOdEejVJeWM9UTdt
T5x+HaD43VwkLA3SPX3ysLjttHZOUoIMrAXt6eYwiWLNNYd5tQ/v2fXsABTq7BtgI4R7KIZe7VvI
GEYnLn//P2LQ5cPL+h1A9Qoa59NbuzTipL1gbNygVmQcAJ1KaQaU2iUf9zyjtFRsgUGqqDvViocs
NQ0vusS3QQTV78lVMnHJZtZ4vNxp621+CAGipf4T+459GfoRdERJXQm0EUsEosJcIF4GEu6OYf2y
ac5G1ThHctx2C5oDWeDqFThFtPA1+othHxpxQL6bpR45vGc2zoxqXqWK0OCOlap0R0HZEfKYAhGa
5ZuXReNOoiz/OV4ATGKfY3QYwBX72Swe3NUZ5Yjy+3tzpRFSouHTTKlQ+sOWyTsUqrQUl0DE+GdJ
JALja5Xn3oaBSE+RVK9zDPKD5Tvtw948o5f7DsUG2KAtOrKG7CKIl49ocbg6kd+wPPF1OSJkQmum
0xBNT2T6RgtzRPAI2RNwR0Suv3r0PbWEab7dNaeJIfZwUEYSmNNtdRdxXP6tHcJGMX6Xj1JCId3T
IwB9qLUkbmHgzt4vme90fQKqlmoxPzcsNqzie5s1rlS/IwRedpWJd4/5y6DBiJ8Jy0GFTjdDtvkJ
NDWxBqkAsD4BdA1w/CO6ZtFeigDB6pXm1CYokplenp9gL1T+VWUAqx9mgu1HfJw7Js6/+jYfb1QD
rLfda02n5qQvfYjWZyJaa2cVlNnlEnxSJjdegr+QuhphDO4UU97j0zgPSG2L7iNShWOQk1Aywmxx
EFsOrTEmwu812f8xBbeCQgdTzmAy8RNoI5dRcZ+2XG419lfErXTNem8g8MLiRh5IIN7OzWmrmrEw
M2RrKrturoBAUaVc9OXu+QneXgzW/JrpEGW7ifetv3lWSBEWxBMKibo8QFyhcawWW3YS7zNwgt+A
+52DMsnJ29Xr4tXh6sihf+qlMlcbKaVjcuCVy47qA5KPQ8A/DSMGwdAypvwVYF5V1tkI00JwBO3J
q1V04YEZ0oV6RUJPMB2hwVcXp9egfj89zUNdKXsK12OC1FmKQK80DxG0/CCeT1UZBHMzwQo9iGns
+ygCt9qEC5izCd5i9cfnIysYG4iHGTOmncVsyaXVhbHSQibLcLnoskd5p4EcbnbS1ZNqF+FcPbwR
zFw8bqwpk7JbSsbcObKiarcSczMokS+ODLjBo4HZ9OMt/gBtDpG9fiX70K4mxBH7ZonFgrM2M44U
6zPk8msgLbmJO29hEj74BjyifmFqVD2iG/muM3XQMZjocuX4Qi1BCc9jOfYZ9i+p5+ZEOVnCTAuR
mTO/r6tjbBFy3iHaGbmK14sNGuSlyC7vGkTjUHH3Rf2sHJYzwPMwweFAn6cN4NOHLEc38Q2NaqCz
Z/9JGFEos8jWnDuRz8+obKZO3Y9/rCGFWRc0kelaHl/BYjZzdVAXMANpsIiwADIQgqeDFY/d5AKd
pvp+uQXkdWCnoNzC22UXQha6anUg9SjZM9w3eJsR4R0BUYPypX7rUpclVq1mJVKtlAyrR3pwHGSO
HBjHPFv42GU02w4z1N/aKLLie2kAs+may/2GXltZQ7rE2954+15cu9SomRju14Q9kxW55g0X4nw1
zaUg/betKPRC2RsD4DpDe/OJjcPw8YZMq2CBu9aUIO94s/+0P2mT+XbRof9PrHu+EYg1dOggzzfH
LrALKPxJd/JLcgfwPHAshvmmEpu8ud70PNXv9IqxwnfhxAoHiioRT7vOM87U8iy+R6UoBfBZEN7g
scj2VgPrbGYdGBm3l/UDmAOoXG/dLDlWfPnoDhKFnPKQNiGvLQHeZwJYH2saTuSqHjnH4sI5E4oo
2O/mSHfDmYxirIACI1gHPD5F+/QzZb3lX2668WOH2BfhZJSxqz3nKlsqzz4ee3jfYx7JDKZpt+gn
ofpiJJFrplSBdxQhQN+9CKuxAtqrvlYPNBaGZLmUs5YKceyc+7F5K5a6xfc5l5XkEuBG6sMLy3Nu
AtnaEf4rHL9Tj1M+pAXmHvzjF2Yj7KaCKrTYLXy7+RlyBj/Mja9qJXOxU0MRlB2KJHfN5gQCaJDG
Vi5+SW22HpdytSj59l7wpaNh0IRq3uuKuhoZaDlnIM4lZ0huSWerL+I35GvpeeN7D2H0OYhCd2Un
I9wGoYL/1aZxBheFZCmsEJsZfTonAAiX3dJgIr4mOG/0GLoRNNVHqyhphsc11Z49Frj0d1DSk3Cc
K3a2uXg+kng6V3vrSJQ7y7nKFUgGXIV+pts3eCDT/Ve2MLEbpTXLsYoIs+zGenu1/41Kf+7kgygw
wcbY+DkeccgsKKPsRvQB+vPk54MU+RKqYjLYyNEs0K4HWbkqhx60gnxAHosVHDusQKbHKsw4DpVi
kaWZO8vXlH8V0+pnpdyFyim6jfm2OgGoZJL18DkPf/5R3XQxXuT3b/rxkrCWTI0YdcgVdE6w9Sgv
AbF3s07duoSUh4KZqngqli7Y5Wk9Gtv72Aa39+M6rG1dRzdX8HehSbO4W0dLpcsS/wMHx3aqtN+p
ruFb6AgzXlzEVZRj2LSq7gRSAsFm+pU4PN24ys7RewWvlOi1pI4Ye/DNsblUK1mWa8MjQHLo9NuN
pjIEegYTpIW8YSYaIdIomsh35kaPJTZcCQUj1QeSEl3xX66o1oAT7csFdUo+eS6L4kgXWdjvFR99
xIvXlFvkGjw+1Kz2Zym6qwx/G65u31A0Uip4ECQzuTuubSp9pyv3Zz6kUAuRDd36moqnCJX006A2
zDwzdPVX2aCHcrW/j47s8ZE5pWnRvRRX4CuciG61B8EG4gxYFEavWHN2tF3rRmuDdDC0pZN2yd+x
mXtbO+g6m3PapVkTd1xrebT77HDmSJVgavJ01XmlBQhwB/xfeiAWtL1WdeoRgFBE02q8WgTGqDe3
NtMTp+nxKSXCxNJXQ3SoU5n+NJHpOeSofNgJ5P8RkqBBLZFRrzB10r68VktR56N+XPHDaQJH8GY/
qGuXW6Z8ZxVPuXzjnfaNgRGSiNyTUmRLPttBwpZYPB2uBk4O5oFqb6LCO7Y9/2bANbcodFPhlTv/
vzw3PzoV/ukUPPhXAnzOulS7iJD3gAqXj+3MWfUe54kibD2+iB1sy41M++maFpH1tzoWu5U/fpHn
s3/8fPYKbLHOOEEhxkgXl4iR4fKm+ANAxjkj79K4atmUyQSShh1ggIDeiH1aRxg5l6y9flE2V1Ix
YqABXCNcmfBnzjj3M7BKIT5cFd0gyHe0/T1/MEeUYRw8EL3P9cuHK/PcZISPEDsSCUW1uOUFgTF5
ofc7L0JJq631xBucoIzedQOD4f9LOZ3yUNkc4Bky6HQN6Fzv1X0QRYAreKKM+XmUOE3I8SI5/zRD
0rn1+qnGb4fwBefCVZoKX5aPcbBRWvkuxQJW+Kt6+zIdEtL+67J+BJXnKojmGM3TfSkHI9VYDSHT
79DV+9orvm4KMgFYTx/nxVvOELyPB2chr0hhjya8d27MZGukj7fnYyCdxgeNN4usqAuyqqugTTDF
lUzVeDRVZ7hscCf5J17HmfeY9Af486nA5smk5ZbeS3iiMFoI32s6NuCdV3m0+NL08vBAlZ9qAkyC
wW/Lc8JLOrHvAeiJ/KokSUYCj0JKwevHwXk9rdT3iZyi7b/N5XfhHXSNvzvPZIK7W1q7KMe+QeSA
/jmBk8dgEUqM9qsr25LmNLvKvF4jCOvGBmzi9/22Xmw5LOdus+sBhlIm7OqM00vlz6MkIp/ksYZT
fWp9WZxEKWLCk9G81Jty7vasrM/1mb/+jSQlSUXt/TlfBkHE3e3eAFp966FrJ4sga23U/VqZaNNb
be8rnxnVdg0quggnBsJvzfYjxPk/0Nl3nBW+uyyOTq8xncOy2v8ta3rgISXRNV1GkbMUf/V+2XSB
u18PbhhW7lrp0TLnnoOSjiAvL+LoDDKBCTg+/+AJ6RFBVoDF0CvKdAL4fVGbrdTYO9SL/2onVv5h
DMbQiFMwYb9B6sF05v/7rq97myz6tMNrNkH/TCnqIZn+lRYrRNHYfZTV9msxJe/qvGCmLGYeqVz5
0wDiNvDFz8piBNiGkpwQszSLw+KoZF1PQ8i7CsfkwLT5O8BJBgv/FbvxJ8I7e+JUVJTXQvPtdmm6
aGae+Wz+CRYMSdgJJAlSC028ArnvSIThVoVnayUMOIq09MUCVR8A2e8ov3tmuQDOBeOdq+bAVSEJ
ROkcD6cT5vLdZ4MIIvmmeulR+qYEWX1YUY04qrM/mPs40a5e9GPegsWHNYpPd5dlmt/UAeJk9gfv
Du25BHNKc98nUqiznwX16+O9cHsoTfyjFzCjcjPVgyucwpAfMV913QswB8HICyrQmeEJC7UEOkYr
JvRAkgivZ1dBgH2ZY5xoVA4HBD2iZbx2FnlVisrCFvBW5oNNw6H1u/orCXfRyKWAXUtCWCss8pnm
yC1sV3Ijk7SVPdWzZmzcC5xkAj2jRiL+tIuIr083lj4Dk47KDvG+J0q2So48WZvW0ULEOKQK8fp6
nSCv0OSW0mUduIiHIXCZL27IP/0sAMa6B9NtoLcOncr798qJ48UBUrElMa4MYa15Dg9sMnbqaS8p
I4M3IWLPYrqAKxkvmu/npAY/gmHtmeOwR0BJp0wP1LK3SLsPps0TKwpa2nf1Kn9QnDBbolIXbK3X
NUyfINJROLt/szQ1EOTa2wHLsMjzTxPYRIaYvPDoL0lj7lFahmKOh3Fx31q0jT3Plf2o8Me8gyF9
Up7soi547y/s2dEZqLpqS486vHfELq1fYISHpfKJot0GzhNEnNLDWK4O9EmPQ9iEoNEshg9wEx9+
TY0EZ9FuUh4LtgjZjMMtZtFWMBtwyYhch2IZ2DEb5YqDCNjQg6lewzo70pCsRT2I0WlaAogXxCig
rMj/bkxWA7igjjO6ko1I8OK6lnS2itBtnG3vtQdg+wDof0Mt4R86yvI+pCuCl5PnrXVG47gAjR35
badodm8+SxWDGsl6kk5ObheynVP+T7xzeCigDQi3Za5pQThgNxJ8lRj2xurgSwczCurizW3VN34W
C9uYwlo+KKLjueLFbHbtD6VixhGswDruEA+F6Xt6u9n+wKssyJ1ejchTy3naHhlrPFDO4mO3EJU5
kO/ZGtWcEDLjvpKh6Uxui3QuLQJ/B8gLNdWPhhpb3ooHz/ADJyTxxCzThTMRmHUlUqGqWqw6u56t
GBGRtpSmZ6rVzEhA2ZiQ5Jxd7jNtu4b+Nwx4kaNFHGMiOvTsNu3Q8JeXay1YqixRnVH6GtdSeHFD
gi/0t0mAHjgZjuPQK888RreaUjilm1PMrS1S974E62WJr+tiws83LTn4JV5qZOESk96rclsBx6Ro
I6ORKD882b5qMPJqOGe4LVd9AYRXNj1NuEMfOnDEoj4L0nRmAudlc/XKJ6vmwGscAZTPjXRYI163
wEWDlP+c2d9Nd0WAKj3kMkoKHxOYHGFqSw6G6dHfpn/nDb7YgPFv3AIt1zUI+hRJ67fZ5drd1cDm
vZUgRh3KxEdb4GdB855aJySIk+iCinyRca9lMZksgW5JBvClWQqTartVzvRV0eDnxvQqnmw1OCRD
ORmerCr21HBrPspET4b3vM35nxGkmIdQAKVSrnw8agZaZHFSAbm84W7guOiwtZHBS8VKca2mhDZ5
zlFwiSsbzqW/zSDkS245JlNuFmkOpYIZnioL6diXNjrmiSkpEZm3/V9VwbehqDVY/tBKpdXua5ME
HjhGXzvSpCwXSD+W9+lyf/hW4P0y4Mocj1ko9Ppi6UpSvBuiv2nHahMZqVAf4XQ7XJCvXlPUlCSR
9j58b+G2fWIgX0gdSCvwgCJE6dyxn1tSosZ6TnwUMS5MD8/NO8FtfF4TTuzLtcW/30t6uUnDTHg8
6Sj12TqNJTG4d0DYdDJE/+O3gosbn750f/ndPzGQ5qcneztNBmzjxccfStmBk+yw/mcy7hizPHp4
+CFVIPgN4t9Z4vb+0ZOVGIDZvfDVEoOY5MM3hSa6xADDTBKo9DtAN6SSgeNRKEgJLATWdFhHDioB
6yf9AJqfEmHmCfv10G0u+IOjhlPHmGfrGDCMoF5xjgjUc3jcWKbL2Fw0ECkcCowaLMMtHQ0Rhkbg
1rslF+oZAnraXeL3jJNO76RLPZAl27+xHvg/GRnBQdBbZVcCWTCUV/0iB1Vxo0sbLz4SFoYVFJDi
RzrWF6rmbky6dKKmJuHKvy3YOnXpFPh8DwYlSvlC3uxcW/uq2JMnTBjENeUOUMGb3wN6Fzah3j4h
5dVTNpibdRG0pFBJtjPcDqdlGD4L5ELNED/Ws1smhCCc6IhQgbuA/ZX/QDLrn27V6TpXIWHpZka2
QShSD70n55SrzvOhfY1QkUmbRxyWCElNm2m2or3MzspFXU9gA2oX0QvHEVWztfYpthQlQMVsE28u
xBXZuF1E/xGYQdHUv+gPlIsTsbtmJ1ykFagNSvwJJ42YDhdX4XlZ/bCoYM2tOMyjDXpvCtv02J2N
3i5o5q7lGtV0EUpqodyPE+wUxgErUrKUt9OCAd+dTQD9bO6BHyvz/PcKSAbNfrjHoRAk3AmN2Q7h
IBPDQcdbE7NghH4T6uW4JNUyNXtOfaY9AyZHfnrAwYNolhtRgNa64lR5L8lZI24TAAELQ/ehVJEB
kMnrTMJAXstLguwm8ESkb6/tbHi+GhmzaGkqrKvcHjiqD2ZCL3igbywGr2sJO+EaoHsJ2wp2r8fb
I8DJtc70JKyCTiVDXbj3GmvWv6P5p22dw8p0AGZWFR7C4dWTjgIvJvOWdbFY9pHNjU3I4ypEGO4+
9LWMX4DVJ8MJwaktxJuZ5icdpBUDcByCQr1JjX4Bn/9/+P9wx7QYCCk9vxwnwPOMFIypnk6RlTSw
F+ccw2NLGp/eMsscV/7FOPxyAFrC3u6yoPqaRxgpjKcGeN4Gcowmd6PhIRBOSILe5gXxhe94sr0p
wR7nqt1tlzR8k2Q2v93NOYzJqKj8pg9uShi11avwTNm+uYydWTRFqONROTc8Wn8OQcbyhj5B9GD1
gO4Do3InDa7zVcNeSTG08sxgmAxuQFFPiHRh7YqqHH1KWAtnniAp0j3+wedcJpy/8jTtOV+2vf0O
Lq/FKfEPC/9spSOJc3IeuzB85wp4AioUI/WjVSAIDo50OYCvr+9caKRGR/eYiXBOGauThualShRt
EPI7ORtZS0s5MbL7dN/ak4wEZCdj55MQmQ9uzMno7GnxGQV+sdOh2spSYbI4jHNV0DfwavdaWo2K
N3qR6pR9zkf9UAbtQgG7Q2G6YJooz2T9MjNo2YR6dWOXBwIeSEVWivPeDALuFiVAE9YwYyBbBpMU
JWDlkMQToVJ4dh0XNAqedCaPNosaPkRuLoCEqsyeq5Zzd5zuFPiaxKSNvc00E5616bmswxiC+N7s
Z+/vfZznto34UVP1ddCJrWb8+TivjWh0ZCYXlqfRtIKttyyEhiBBo2HNW2P+NUFq+RiOIuaUjqMn
bfZ3e1RPaCEPPyYwcaFGEFTCwYaX3qDa3HNXpaWXV6CPXOHITv+BFEFK1DTnug3hYGQ1bUyZJD5F
4OXj5P6aVVxh8NmvcJBNrmyqwefQHwmYJMpKtbvKdGBQcdOKqvudE4Mm70XUMX08lwRzfYxzkxqy
5/WYo2Axqtt3BclludPNQ1ZZ/+nYfJXbRH+AUXEFEMfDPzB16dAdaDU5toifjAdcD/pEfGY7fK6g
c6Bv2Y3CoVBkEk7qC5/kzsYwMiRXHZ4cBFOqX0+kiNiHxvyak2zQzNGBmIqYaAhF0Zh+XdAwaaCr
ITQmCMdQmItsgjvFI5kVMGJcR/3lg0m87sm9BRQlHXhI5kIGf6jRnLG4LG6fdW5wBZiAYBmBEQIw
ok9+SiLHFN7OIm8HCPH8LfFPuCBt5DgacROkpIUduM3qY5gptEy8blFl4FMpCD6qz65/ut0nwXiD
x4gWYCpIjxnmAHP5IYoeKc8Q/kJOb82QqsDZXr9cHGS31pzUxMjMgOfiw781iQ0K/ynzOQVVrNXq
GuPEIzW+IM6do6FW4/YmpHAIZoxOU/xW1Fmph7v/oJtRB8F8ZNS5XjXbWcXktEHOust3CO3fAj3s
OI7dFfHEXIOIqYjCwvRvkqSF/s4msVj2WEk5zoDUU/8HuiDZT8zkT7Po0V+L0kAYdkMhKwxTQw/b
zePRNQNiuIiu6ucVDzPGDZ6uurJcYA8Kmis7di2CuSPwtVUq2bIW4VnpUV52qUdR8zcauAv+ag8L
gzWDyLvRzZVwiQi16cI2LrE3QGyB68EJxCfJMLHbie5iJ5J/Efpm5GRkb3H1C5XeWCyKyECHkDFB
QJdcwzFjGgZiUiYmKIqi7rmyFTQatA8DGWsXYPt/c3hCh6Q4JU0Ltootm0yKoePvBJIhp7+aZT3r
88FAc7p73uJreyjDOBvYdgF5/2tioTqlR16KTN57DmH5ndieNSdarfsXIaS7VyVEiYciFlonSX9x
xI/IsrbzJc5KcudylAiH9+1tuA4PZuLGZoZkn0vwaBldgpofMofD2asHGhIYQB7ktgqTU0AajArx
dAvvgs55WEaACP+6LqXPgVnIUund0bj4kY2a83Efiia+4IThBiB+3QObUWT38GmTLpgIcyD/eGxB
LINAPT2ffqtRsgCAGXWYiB3dJJm+E5gs0s/mZMbCzWY7XGq30Ijydl/odULOrCf+BJnoPW0o+OVD
M42QzmtLlkhKN43IYKlNSj7hvNuAcRBh8da2FgQdEC+Rw6NhjNXOSWNMl7yP4zsthlRW3cco4gCT
l5utWwQvlWBgXT9WRzM3kthB7WHxDgAlgAr16RmdZYZndOXsEewMfH48vWkXoHOQKwaRGzkVhpGK
sGwQbvBKiUAZxlAeL4xc+anCGZIsDvsJa7jZAjuv0V33UH0ftKxPKApujwAywevLO50vKWUoC5VR
/luKz8cBPAmLYWNMLOKdgjSAyTZFTnFVbJBYGCf2ZiAhnYvlPGh1xW21Vf77q44/+1lB5kIsfyZ8
P+gr6c4c1+PdnUouaoSphshTRVpeGZoRDhfwdkpjIlOYURwnYtAE84C4SsS1zJjPYDiLy+OTIf4p
9EkA2BI3lImgCi8Ucvv2l71upFusKwN0jom1CIPKWl3Tvro6fjquX2UXTnMEPIQlLT/DJYCkcq3B
TkquvnQ/4nPl3QlLtz7sZtNSYEDPFc585HmzNI/WiuuOam1yrEHIy7cHjbIVREx9Z9Gd+qB89IXF
/AHYs1GdJBki89ZQXAVoq9n6z3//Rvl70LEBE19Mf9Oa5jN2A8mAaOQMnbtC1zOxYfIe9JlbhMys
3Qsy+oanbWVvUFYSMKtzKUAVlKP5/DcQWSX12jyRLyLlRkY1sQ3kiUB6TLXrSaeaHeBcpWOyLrZ1
2JCzs73lOldosRQRCxbWkocaPP7YOoPRkv2S3ef0Lmj4/uOVeWCPZDZUkgtcvilRIwD6E/DPiQxp
rZWf/W2UCm/riMCFVX1B+5uAaVhNtCkaAYdkMhRHBhaEokmcnC8ZKtKz9uQyBdujEEN2HZFZBZQt
yVdntb/DQQUB9rFdQ6wiOF7gZEiwap7u0gwq+Gv7NuedXvHm2zwuLWJBcSApZ3Tq9J0652ZnhmO7
pOvzrk5u+xsWG53BdtVavib0Q6WNVvyoWozpM28ONxBFRMuXFgEbKKUjflHcG+bMrWG45mNs5f/B
P9r7Mh4NaJYEixhsT8Z4Pz9vMrwpAk5R6aitj+3BYvYmmExqOlFC/Virff1K0irfrKAeEiIJ87sJ
FVqoZnKFndxJcmKTw0M+NJFoZuzAYKII7a2pjIO29xXiS77kLxyfmJx3wGtw2sl9dpbNtgmmKBaI
zvBZvZ2zfK8NVs+GeW7/u8gLRA9ig1RbikVAntft4FwlxQJ/jr42z5YQwamlEeJuM2+n3xaegCFT
kVUEEBnrROY+E8kJO6tT6btC2+jSI1Klo7xVY4urHgEWEly/mamlHLp8gomXEa0IzIKuyuhKpXPO
YI4jdn2lRYuUqaUfPK2CdylDUxlZpUqoZ3IopyxM/qu9dVnZCVUxgdNKmNV756VbxjSzWc6VRyNe
kBfaDrDGgOVJ7jNSseBMkt1lG+c0oWeLczUeTWw0cbfJANl0GZHxkA6eeVLakxvIU1QYLfU08MIU
TaLl8K3XOU2SFAZ+R77SDFaAes8zkbncjoP6X6Cgu0f8GneCPDYl1Dp9XZ+JMQ8VDBmLMWeQEQmw
EDdzNzq/B+tJV54a3hdS7B/QSzXDABld0yk5hS5AklrEDO5M6GxABsmCPK+G8aoHT0UHip1W/lZP
1OJPzfO/6ZNZN71o6Ww+7vZlwMRr5P2LNkboUqjIYkDHMecEuJmehfZmApaqF54xDhdUpYJCq1jk
ybzXFVLY0WDJqX7oMXg9wKMdCebmuZmePT6zG2AEz/WO9ajnp5gcD3aqiDstO79hsN0Xv/T3H0As
qCF1c60C/g4kYG/B6u6DNRymRUVqrMLAikr0jhamVWkM86EK5KnSsiR0caXXG6rN1PyJzmqH0DJ3
4LuigbynGfGtlx7YNTuKr8XeVVyRhNKUB8/CT96QbomwRTbEdE4vJh3iRVqeXGSZhZUAIg4gBAmt
HcXr08ViU0GIa4LEazyOht3AlNKu6+rCR3+24o9mqHoflleFgJmnE4EDz8u0Jdw4Tu2tQDihOn/3
K1JFa7yo6wE1Bs2ZyemXmnPqrlIKDoh07nOGGJOav7h+SPCC4RG7dXYn/4TPlNQGrTU5Ii1KLfw9
bKQV3dXeupLB/OnlIYzbgOVFnFsHZJBmq39riQmJ6TSEPB6LqsTHbQ6DzweAXecUUSuUKl8v20et
99+isHpH/Ck7pqUI0WS/Ml2mMiNZEaZmZi9B+F/HbYapBK+O4dRUt0zdMEBExF7hzqmITDuSQhOQ
prsqiKsBJIK7Zi4JpcJ36VfhIN/bxK5u+hhi5y1GAl+AK4DWfAjf4k9TDypNhb2l6xs03huHi26U
yWaM3FJURKFK/pVstg/8YFSDfyZbiZwFX6fy4GBp2WiyL5WGeRKegb8CtnvqgGiP+xuBu92CU73z
UZ/6IseHQKU4BHBhpzTSLzm/ogHWjp7XIeFZdDf6RiOyi9xthcyY3STg4CeS6zm1xQHyJVa52UZy
DP5xLe8sqzvW8UiRMHmfYbNPklbUYUjdMConRk9P7t04HNT82DB0hRlaU3UtEyxOvZmuF3o4Ex2g
oBraNv0QHPVPU7o4MGUX1LYjdyQ8650Qc85YBdEpqpBkAOrjFqFLqLZFj81AQEUTsH4PlwPU07R3
Yn+UdgpVkV6zWE5UdB+G2fKLWJgRn6pWc0zwuxRDeaF7J+dDO3LNbOQcz71xOxaziD4x4hH3GJDk
+U0JOsPc+ptkAedp2t63e6yDQzrpUXcsRT5XKijvc89Ud3DlNKeg0Xy2EOgcw6QMm1tWATzqgo/O
3AUJUb0f6cZg94j4LPemnt3k81ZiYfU8L1i4SY8d3q/KeDmqV01FmgA57NlJOza0Ob/iagcmemDX
f2Q0gEuGbiJkzLKCawfthXX8t0I+GBqNB2kuuQyXMdSyP2aQMuz1TEl+XC4mWsQ0asPe5CyoFhyj
51+KjarGrQmIw6CP3tcVwxKmngPzIy5TnjWNcF2fY+NFiZRImzNIVCEbCcc8vkz6QK8Bf2QfP6IK
v+E7q2kVrqsP1zp0z0SyG7gQ2WIomXyWq1pLz6rZs3R36BfC5zuvkRCWOL7ShrHSYrg2ACaDTYcs
D0eKgV4/5JFord5vvZM97bsa9SP/zlIgGtVDL0bkFdKcZKiCtoTBYxN2VTYuxVjUhT+230evDu2K
fJPMujrUeY2gnVkBfYZ2uEnxxofogE/RKUJW62pM3PIUoK0WLmxleBI0D5qQlzRDkP7OFf30hwyI
7MfgV74JqUPQISenCaHz5NrXeiAljMZjHd+ewRB4QdR+CvY9q7T6rl/spq41WdYGbFwAxi4cjLm6
1wt/RYh7ehtt/01SO5jhEqbg5nAb1Zr1dcGbiAfeKYrLZcRnvMtdeFqis4k4bu6KslvM806khOQs
9fkj56nLZH0LTInG9LQEMuyiuawuPd9v7n6oC+xLFZdCNiBo6BIyswQEFIDWzLuu6EdHGc2q2Hqs
loM18Zv2py4Q9nrp+/MrMMyc37sPD1AVA7n0Hv1mf2SwtQbMVphWbz3CyzD08HBdRLT/lVKNqVZ+
zGEywNhKd0wLkkqTJHPOjNmIVgkuTwtBw70SUJnAhhZ5GhzxZEyKwDgjhevCPAm7EWnNNKCjuUD2
ybU6qX6OlJ/MsyQYjqq1A5W6ii74PglTgkIoaPS/CnKC9XMJBHdT1VpeIoDNgU2LqJeWUgZBdJx6
/b/e5Xv65PjvfrA8y2OD5OL0pHqdFFND7ET7PD/rcqYt9q11X6ELlkRWHSAQyHUO4h1EvIoXq4fx
ItxsJokg5gbFEeU4Bo+QxHKxcBmtT3k+ViHDLahm354InKysDyOpdoG8F5EH0o1fejPlDBNIWSye
wylldXywwrojhgIgTPcu4RDu/EfDGXyilNpwfF0IUrzKE7Q7Zr/GuVmDvSg+1AwmmqQtAeN0Qeh6
nqNAdRExqE8soEWBWNOKOt4/gS7HRgbg7ndoFhke8mGm+ICV6aGpaBs8jivUWDdxoUsHdZJfzdHv
HfGzMaeA7KJ2TCgJgQdAeomH/GmLBC08FKQ6juWoP0Qu65aQB8Wvbunu3Jbf3piL/mnC3e/Da5hX
fD6J316FG6zUM2OzGrO6lT7Vo3WguY7Tra5dbRL7rutPCcLx/537tCXyXkS8qh+U4J9Evm6IZknG
uJPb0XepPBobr0QYoro+4yCJB1aDVs3fIBYpojuM/l6ebAdELEbtH1d7Jp+gqt7ZYDJMMXNLQEna
WlDrU8w/J5yBLzMlbHtdmXy9z7BJY31HzLCeY8ANZbSxjjRau58Q0mLSsQy4zTWq711OJS0nJPyn
tIAVR/N5kGjC06wOHymXJZzb5+nxv0jstDUVts9ScCLmHIlGD389nY454+VdX4QRjoPeWYvuKefQ
2c6vLZ2HFaosW5vuYM212zgmSwM7yWX7RRbIR6AkoTDpQKUaE26g+HFLaK1HEFiF7My9W9krXBFd
xdx/m1IcunDQi7UVyn3ncU5tobh9XrMak0mrc+erDkSu0hQxMfAZsFz2/qUvhfqsFTRUj37CgpjB
n5NE5NRB8gICWUus3vIOwdUmeSY8vKxs5FdcgjMxBoZ85hZOvuDoavZslrldWcNClKhMSJ+mS3lL
UscOU2rFHGmJ/Ib/Err3YhY/XVQ67lxAgBLz7FdF1c1x/FKX5tv2AFParFELRYZipCUMyly/X+Z3
EvfKj/D7g8Bx7ntL3yCp/T4oQw2IJ+QkV/DRotpJK0dI3mYGXvjzSFl6+8oYqFchbFcMYDfUSOas
ImCN/E7CH+jVk0F5Jjo06GzB9WgMirkQ3Lx/Kfyl5PKiNQY/eVE0INxh9gsC34oBV4lbyq4ZmyAw
1IH4YBgCMOxrOgxkifsORIka/anfzWGUmDFNkTDWUxOnlAcGQDk0OIJw9saPXxkzcPbpYaqZiSXv
5NEwO7kVRou+fco0UgIT4pnd33E3Q94APT9xfVk7POUt/bzbH/SGsDdtVvYUKvtLf5WBx38OQd6g
AmR6K4WDDUMlqmUKnUR87rXyFPp3Be/AHc0PQtMMRJEAAr38cC0ZSp/G9gh2ugQXbnLaMF6W1pcl
ScSPJZEBzTiZN47nxY/fnHLXgsLzucL4jCuCXgOnPlpyoGqA/xqx9vXaifqIDxJnC5aR7hNtAr5K
rxEJDgBC4jXLORtgRt+bBBonCJKqcwBbjYmd9yidWxh07QJtPT1/eJKVgxAB5fRV+Adk8xGsz6c9
kDMu4yKRr+khhZiSv+Y9uT0rLwJGAq8u9bnUKisZwAUz4lXRkp366tGb222kjR/RDx+0sOHFhR3B
LOQltzTzoUjacvnnELcpVnNxIaU9r6OcfYbenEoqcrVBFN71A1sQKlRozuVgpRU0ypAA5ObSI8/I
OfzZ7VEEDr0WGSID3513CQ5ma7irRYREkEI6v1/XpoHH74AnP1tjF6lApsZ6wLlpXOBgXruUYXRS
xQW7Bpoa3xV9V9UgZ25/2V2kq6Cqts/8FdtWpHACHoFiwoPglhepa+MBnJlssxovCQ1VaffuAj6H
gPY72NGsZw76amRvG3EsSlGoSJ/NbY5QIZ4JajRwV0tzFJjJ2CO3IwFM9TOb9RsPvr+o/C0xlUG7
pN7p2e7qKCgJZIA6oW4okd1nadR8oBh4X7RsqjJZ8fFbaBSkSKcXcwkv4VLOLjXmn9rFj4o91ouQ
hAod+lKSJnR9e0UWWshNemipXehll1l8oIZeZR5oC/L9FzYFeXg9bBL8b0/BRb5K6gd3vbxD1xWb
Ep2q5ujdqXHLnp3hADDDgZlHJ8VEZHGytsiZKhy+OPI9s4RRGPgJrAoRrANU6PBMUeuLge8L3rRr
rpIocci7XYnM+VOVrZClmc9uuAxqV//iQxSk3yURlR4wXE67Xbi66TU0dQpbomnoivvx2QuDbpdJ
NsBRj1qzHROh3uP83Y6jAOEiYtAIwp6SBG1CeBnDvNTJ4N0tmebgrfrSXEtXL2iNJNuS2lidOt6K
G0rOvR36LifoIlkf4QSbzWB6ArFo5YAa4BxJeICPmXfEMRw7Am8RYWi9hwnePi6+QcE7gaQsOH9g
k+K0zSArSfveDE0xhLE3HmbsssQfA8jUDzBSOCEicV4Y5ddDpyHS9HwtLSppZnRImG4oQOz5ZSCM
Fq+5TUgLgxRZBsle+GIW2KFrqhS4d91RiQTwAix8taMs7KVyLLFvrMc0citKz36W5Zl5YGWloHbZ
4HuXMfnGpu66BYZd2FYH+c5FV5I8j51Bs7eW028EcKIhi/BwECgUpS4fSLim1F7+YgXKZzoGqw2A
/x6HT90T0glxzIeG0KY0WO2bjRoTRciuzOX/NIw+M2svLTWe+mo+ACFNVL6r4YGlOLNUpZNs9mst
MX8exv57ADn/QRceJpvXhuP6q9HgxIxE29GQ7uWtNZMZIqSsGviLdr54NF1eXu+2+82pdvpIx64J
tK7/617H2OGQsChvAta5zllAnNBkojEoyTJ/Sag1mNsRh9HgXWgRZQ2kD91rUddwP2NWB5P9FyBb
pj6flKAnpry9nj7UD/vPwi+2PxHC9Fs6wYvSF3ULlOlG2Po8hFZaXr+FL5QZXwaBgCJ/qWLkCPLD
kR76wOGgbWttl0byPo4eUw4N8xGHCgjtMonWYzU7wwpovwiHQAGxAr5CZt6L3UAaOuueKUa/1Js7
XrqG5dL4CqxpfEo1MJrFJiQybQykUZPZB9cbyE/6LZ7ew5svrcT3IYyoLYhkVBNoyGwcrctnYMlu
xmVNLt378V9AF4xrV+CJ65ZDmVWkDSmLs39Xpmk5c6kRNwJXvIZ7vEHFu6AbfFqqKY0ZuBRjZUvp
lwP5ZwCg8Gcbc8QB6ArRwPbFXqxPvbJPV3H6/P1ZWps6t1YUrFwgDLFOq+sBT6sWY/glhm2Tl1Il
PAao+cgzJ74gZtPuHCGV878SE7bmPQjx7tPmsE401Jv2GsNRND5+bDNUYfGeyswkOFZXpZW9b/rK
Vfe9qUBe5O2uYyTSFTIsztBUxSxJLkz3yHxC1Q+Y4VUmdiHoLC1CmBhZD9yzxTHfQyyYmDti6MPe
b1vQVUpmN4cEXL0URNd+3PhGRmcn2ABJrGgxrjUD3hNeAwttlRMQJWFAPpz5mgZaVfDhkL7DGtdN
y0ctJn+hpp5P7LHR3nn1j0GdipHf/yTMT+wQZcTe614/H6iAgeTFb5xYHYkn34DdjXEav/Xjopow
rS/cQZw/ajwzInOCK21ze02+d2V9D4hIih1NwlaRSTGOxUjEN+UrwTHE4YaTKrYq+47dboxcgLmP
Wz1Cq1ISKD3LBRrIJAIcUOB4hGhWFOiJznttaOxKk8w/2y1djMoeFLAR2P5G6z0w5fViy91rNZ0Y
Cr0BLHHAVySTN3bJwgTCnA4WyYKnB+DgiCXL4+0rzsLX06GPePB8dSMdt5rzNBpbQAvdIqZXblQ/
buXVeYCQv+8FVkSbCkG2SBoyunehakFvu4ctCgBgxC87U8xWjSXaSYVgMk1DYEU9mgnkUShP6fr/
ZVYtx0KksdE202rUz12SLU302bLaUF8LynIikEm9VND+NjvG46EXR1iEV2w6W6sTC6GBVgFsMayb
hpOa2dA2wOkTx+RY7lkMoSVqOvlcgKuO0wa41uyILvCMv9BzBzQpxpiHR11vhA39f76UhWw9zWh+
e0fsN6SG3lWurbzZs0nXQYUZufz2odMLRjny8p9FmrP1dlJvFytBTUuBHZ83mK+sa6Ybjnpk6VZD
VWUE3hyra+hpMoPSKQu6iDeCiLvOq3Q5VqVTc/ovrLRqMb5HNQPxTNJ4f8GhG1EI2HxsOb6ThS4b
ZFtp9nAgh8qzJBmZ06jSMRqW9p4FocFv8YzKtQDx3T3vZZqdv0weCMnx3vYX8eWW5xZe/iBD8Sai
rPo0ffq/dqv3jh1nx7BDtq1PjpnY1JyRQQvkEUx0wm/55lzHpmDYHD73xsVaBQ1+m5Qf+hk54bPg
JDmqirjp+IKiagsfDtvsVXFdvh5cHtgO3chcUJ49eCZXlwqOZicuvRkS7ReomRGqHMqpw2yb+GXz
yM+KMpv/Dt0tYxWos29RlGJfglI55KYFPE/H/87X9DCEj3R+mmXUZb5ftgtFZ6WGUj/e48XNAg5A
DfP8nnx2RdyxuvwspgtccO5TBep1rtMtrrDwNHSx3EgidAPE8FYTu/7NSwCpgLfw87516gBaTnrk
eNedndEk1+mh8fhN+o07jtewhNIK6t8pslRz3Us9dxUkrMlAsv+PdJD1pqJnvNfCv+ye3hAWchSO
2Z3QJZDGcpvdLDSHfHUAjliUHMHSHaxo9n2F+Tj33l9TZPj9qDUei4VbH7HCyzM16wUBdsm1uQug
VrZj0oVs7/RtEP2lC5oQlbwdjxlL0rZ5CbNE1bXxxnHrGid/zJUsAzcY2pyomrr8x+VzGHEGv8Ml
/D0vZ/h8DsVdd1GtgITRjIjV0QtjmRL1T56s9RlqA9ZN3anenvOS/vDoeVIwKDV66pHgga9GlcIQ
PPdtnNNMURpyNp7FUHBFQLdcnqB2cmSBWEWTz1+pSypilPDrtr5lr/dpRVBl2Zel5SAhPA0WFxkr
JbAIpAvDmprUfK4Iil2241Vvm6N0xvg3DyHljiZqkoJRsWiJ56ChojGL23uDirPd9LRzOX1vxAUF
+JklBmFQNOaPCIQ4FucHmXTqNOWUmPGbtH4HQZzFzooVfgyPf+LvJM/fdk9EenNAzNoFquJkd6tI
t9q2251zEQiu2+JlPpLe+fiip9DX+w1gNEen3mKrJhgx5UdTxvG6YnoQMWadPOIXcS1JX62CBAdH
hFnhWIJ839sBdO73pT/vy/0rKRt/zGx07c/jl7tIcr5Z3eBbTa/cSEBTFHG0T/sdiKqYbub4bzz+
Dn/BKt1fjBxz+KOPQNspv3bnlhE1qa+nyBOr+VroVsFSml9TdOfkM+NO3ytlOx5MJJYfJvHr2DKq
9H6u3EQrS5wOEDbHO4A5zzSWXEtIpOQomUdwhc1cAfNdRlt3yn6H8i26tYz3+JhmBj8EyrwMZG3W
7czL3JVK7wCU7vaUWg4Kzc/wn54PuKbPD6si2+eNlfFa5L1WwRW+ah9AhgoAr7GH6nGAoP/YPsB7
isoImUVWoKc8STa2NuDBBysjSH+3LEjyDbXd22RAwEQMviXNi3k3XaQofMv0BuREky+8Yn/cphCc
ioeFzHNRIWSqpYqw+c3M78kPIMu+eWFuym8zoz3WjIlTrCETENjZ6+qxHbIfUp6yfIEQCwb8figd
e1NU5T2h94E0IHsDQx16CUFHPObn8Qhs7P7bbpdzOI8yaSanvzUfp0SORUKylWk9gT/4fWOsdB8i
9voxSuAIG8QMWfM3ymv0bgS6itDSPvKfjCvfHIFwx85rOpZuquxatNtgYSpctlP+QQkEzvgYErGa
Vxbj+bxxKCMCkTvjRndBpw1AsDnwK+DRKSxtCaBPjRSQSai1MI4nHQOWU2KYgjW5owdDQnTl2MEM
kvw2VslAo1BIIbEGZtiOdf0/M2xaM6m4HJCBTzX6wNUIjStmjEZ3CmdlQsPV8QQkaVTe2o7Pk6Jc
b6cQQT8jBMcnZ21JX9Q5JY95PIK5MOE3nQWxmCBnMJN0rI2+hIpDGZsUvjIJ1Gjc2G6pUU9TC5TH
APJhVANMpSElvIqOc9Th8LB2JGex35wJdWPIvHOqsMLbUosLr6sD8jiepfwZ4wdbeUTp47hF0qeV
DQ2Zy6qqEQbxstR3AsaxGDCzNk6Sk9VocAuVexZtAWX7QSRrQv32Oa5IMXNRuu2xzIZVuJK/GxI+
P67lwMej9RGcjGdXqHmkHUEAaz24FtK2mFnTYGmfXWNY2fjvWp/i6f2eWKTo4QEiCR6l2wBrXKdy
ukKc156pfzXPMWBP0qkcy+7RckXCQUkFoCviHct3At9rwdP/5DpavPmBn+oXIO4klkYiRdjqMcjK
8OZk4TB31bPSFMY6pDbQ1EPvqhSF/d+w6tT+qglJ4JBwDWVBaezljkL7pZ7dyvHdEHmTtwVr+U+Y
rINMSQzrVxrXHMd3lsn976m/Z7PGtg2P81s1Pb/ys63E+PMteu7z6XZyedrY2nmHFICHXsqf2+Sa
Dj+OIXrcPvqesLBASdknPLQuoj6Kge0hpQk8MTD7uy8QRnUYmSJwQ/JHVVDDEfUKdgx0d/+lHMU7
M5vRekLIObsVgIrukYATwEJY6pTrxbQtnhaSuDlmDdDZrt92kciAzf5jAKCGPUh5M9JKu5tSziIf
4uF3IvMU8Yr6nfwKXeD59hoTW+UP00hcayTS6fLe9HmYW3W8i1yquTHjUA1Dq2jrff9+gqgSnWUP
pQuxxSm//ALm6WXvASb7jWsdDa3sJL/ErWByH2KpNErKIdvpIJHDpCQaY5fIEIa8dKeUWmJi0Wp1
Zwlc+pp9u8iUOUdbk05tQ/xh4yxpvUagRLwsg9HGO8cTnbcDDtUosPUTyLUfSnjDQiWZCPq/M0l7
XqF3hmxN31UoCGbUXbVzB5UXnOXy2b7AsbX5H0fHaJ56vnEQnDWsKzOUNc294eA9DuAAhLRlL18k
iXUHrqu8nrNvgbTRfeSq6O2aHiTikgbzA8wfCJX1P/S827S0jb7uCEYMARUnrFF9GWVPjPMjdqsy
djyp2by/a4XtI2g2rKgxpqP6RhghZkYJWor/+ve4az5QnqTltGvsQ+n/PmU1htairlOs7ZUaWRsd
PsRCbk1I4h1CkjYdcMXBwTx5naMiCGLZuqNSWUdwgGVUJ37/DScy5w2G2y8J0UVyhimvRvXUIE8/
wMt4UPk4EWxzO/se/5/BXKouK6/eWqdNeipE77t/IvQ8dakZUABKuiU38XgGwOXEu4YWVY2y+cHb
W8BrnBEuOwb/pcxPeWysWXCMLlwtNzf2bYaaDtzmwL2RS9x2BHGG/qbvEJ0rYrGVF/m8tNpsH3rC
iDmWOxhkMmDqEBFM62nVg5TmhvM5dPHJz52Ar5VfoxlJFE8uHEwzosP+4+JN30gM4Sd1+XUDbrjd
8hSHnUwEqPYx+36Vbb4sUOh3EKSJ7u4jY1HbJhLGsbs5Ck+YLvLu7V0HQu5zdRcPLsy5KazQVHVK
Rt5A+SvOpVuuCRHqsV8ihEbqm+h55G0zXmtrLDwn7gFBt9z4HMTKtv2i/O406mzG+rEy1Rgv2haZ
FquB2dXVsK+DoAJgfq3dJ5yZmlkWzXHIH4lY1hncWCbWOvDYNiMvqkcbIYddwju1hD+A1v2nyfT2
Xdg/h08Zth5LTOuA+k8WiM1PvBYYur2VQlaT0rP8Jkr7GosG1pphZTlUvqVrx51QPcLNnKoG8ope
JxrWdjdIYVz+0p1P3nHstWyqO+xR4W4sjU82AobuuOGLRIRXJi5T1yE4I5wiFF2ZuzJ0XrscBFuW
ySUkPGpANoVnM64pUp1T4BOOzfDLvVOIoDvmmSB9j6IRvkGb/bRxKIVUDaGePcTH65+twmlhAy3v
/dyX3R7O1MlkFhaX8UN2+L2ZeFO5GCXgkm6fJ5kIbBtBnyKJfXT2k1ziIA7hRV7gWd1kUsBZpOFI
XhKEszFx5iMCVhWhnU2ak84yOIxrdmIbZ3RExuolG0jL2YXnHoS1qMKm1GxCfWwKmWD9iiVONLg1
8lg2L8i+uAidrhO2P3SDTL4Yz8C2HBHoUySQqjlZFh6FnP5BclSFU00rdD8WlZ+fra/BPN3C0+Ti
vkmA0zm//FbFJGakkahu+rhZs2mYrS3IsbfQn6GNwSF6nEGvAUFyOS9DjLwPucTHWjRGMbHQS3/4
Do62nDZzfCTfTEK9pyCQYUaMSkc9jrl14DB2NNM2UFozn4IfNMRfwEDbwWRaoAhO8DYsN2SiaYc3
dNCH8V0ve0Q9kcxSWd+aZwH8aQOaOI9r6bLDu4iCewoGEH7BaHGcJHc9BzR94gJ0o7eiBLOFRFQX
U7KKAalLO+/8+R8PwkBsY5bynI90T+CARTPz2jjI1Y0oGhpZyXJyh6gEh866ZVhO9T/wTDKwRpLu
iGMxZkDw1kRv9uXMWyBPrPlQEREFAK31X0vAWaFIMt1WCd/2yePd7NUZljfSGBxnyKRPc/1mJTZq
Pmn5yZGaKwIQelMUeYTz9oR1obT6AKZywzuX6J9yGKysJstzU91MpDzSFtYVpx18nrfrYUtHgEPs
33Lu1oYktjqRbSxI3Q32TxpO4V2DY/Ol71UT6PHNd+bDZB9DwJZOfPJkx3V83FWXypnWmZmzRAJO
YNi04Rkz2wqpOFs2sDMHvZogTCagONCgZZ6o5ZccadjAE3ZDkE0J2rVjDCh02wx9O5aevmVFOear
8O2JT/mCQMDAENLmOcKTIbqdWIkZ5zdkUr3CxPRcHnL73MuapvEDyPS0TBO7KE6e8r8I807oocpY
wW7/FAJFkuPUf/GuF4Cw1LUc+DR60eE3pk0E2bst2YHbpG8qLWabPnEL70LsrXJDB6tt/N5KmuLd
QOxK10zYpJJbsgr+DlHHrXj6sqVWbxqgNPG3FGEvT03hTdSk+ZBgfl1D+M8vlaYQeAtMPrHohYDM
QleNXuVbaSF0O42kd9SDH+IMeWSEDKoUZYbuuS1DSjvqY0VuOexa9iwlNObg17AIjwQIMQfxvXru
pENUjvuBnHXqrFlSirwU213Fd6exX9bQJwlLQ9+KnuAp6rfI+tLAugWMnE7j78cf0uEq63tQ11n9
7TP7MPmG21CsHIXCOCvH6nfcyKB1DmLbCPJCjodJxknyxkud71kwY2qzO06b4mUxRd+y1NCc3QMc
GwCU+lDgpusyTzaW1P4kpsLRIt5utY+2aCDCxKVt+rhj+181aQs2KAvsdy912btgweZZ9kW4gH12
ZeeXCDDNiwMLRHapbnUBdwfa5alynfBcQi6iT4J37CrVlAqYUIdTcWiphWJVWU5aP/TKXyLTrb8u
MZo/pqaNnPpEx6rJEOqcUZGsubvIdKnQKUBvbgvsccmo78ERUBNAX9ZqefmPJ+sdYLBI/BLWptbp
0ty9ZNYvYOtBDurNMvkbY24qOtZ88L9HDoQyXWew4V5hg0QB3I/rsBbIN/FkN1n/Qowg3aXW3XSC
uDeBtffTuNonDmcntCEADT1X2jr+8g/I6WfhUfxX/Iu1wgEM2fFU6bxfxJL8t10cytXqAWAeu4E4
y3rZ5ttg1h7vrndNm/JELoOovRp10kJeSVNqkgSZZvXvFUSx5Z1yAXOFsSn+u62oUZARbudv+u6C
C5xzQZtBU+6dCqruBgLvhix5OZEiRU5mBc6CKn45Nu/9dDXnD9Jp47loeHqYYYDHLwWbgtvxbtUL
x66kyWHRY1YJN0ORL0nxpPF+z/KEkwyQ3pZ5AYt9I1wTQKFCz613gUcbD3VdtLcY0eqRe0xM8xAY
3/WQYjJdKSqmyde0VPt8Eldp4FeS9gpO0TCQGmL8RFQgO2gLrU0J6zk7IgHyYN5MyWdoNY4VmDyg
2iV3w58I42gD6NvzoaadBb16fwkITqPjqQ2cC+ahEMOKVRErI2K7J/YDX1UYKuzC+GznzdGoVibs
jTm+z3d7YIs8z49ORCeIAP5wPYROk8rzXO69it9ZsGSJgcbQZiY215q5YAnVmm88eySbKlR5CAKU
uKEOwudJEBQAQFBpxIWEndy6mDDcu9XLxodEBY2Z9wXKP4uecKGeB5mIKttWxJZspMOxa8/JSsAE
I350cXH0uUfPvdBfa+svieH9YAQk3EBWB0SVNh242v7HYPg7vBVFeVyoNSBgMxJgltgYYdgzpn5t
ZXQCx/Gv8Gsyhyc4Kbd3lim/c+JGDqIldsEo5TRxpmvwoK6IQyGpRwLGXPJYMv/5Jm8IkBMDehNj
U3u21Eg7o2g3s7RInxltUvizSLha0qvpGg/6VM2T9zshsyErmJJl5522TCntPOAMo0ZnN2WnuvoI
acw4RzRputSMBNcJdFmFy3wchrXgNQDaxr18gVvZdJGrhm5uYwWC06vLMnUtwJYz2fuZf0n7DKL6
3FP5ngr9fbK3aJUFsSXIqF4SBBMbtzQpGrtNWWvGNVfufi4BbJ8Yqlh7jYWtOGkP4AgEGM8nZS8b
jiiL0eK0SW3MyHvUJEHEbtstl1C7pA0Za/W3fVltEUxWY9+LeLOK8KPunuyIQJToROTAUnUJq9Zh
TqGlJJqmcEHIak32OiVzNzxxvoiAXTvbh4iEd9dQnKxE+4mHwBC9LwrxQ1YSxTiDd0oS+EamH0Zl
HQWRHeQUC9+ZZXMMmJ+exqDbCVikfXOjSSCFcCoPsh2s2b9nWERkCnMIEvsClrmsQ2rUedyTlWgP
lnC2beSbAed+KQPNNzTUjRIbDIAy1ICnBw4vB7mHg1r42AmWa+d1VTgorcz5za0KKFbyDSL9mC75
2gcWE2Dj65siaXJQJjxRHNZFEWARfGx/o1SSLl+U5yPAVV6nBRAl2lSDZo/SS42NM8gKGo1Rijjm
pBAJvAD4FGaFboql5G/zhv75yNedBQce5BTzmpevaKDivp+8kTNqaMbEPXaro0hp8+VhWIca6Zh7
RgpA8LzZ3pR2stQcm5pu/QyLO5v0Uku5/lNcEkK+LkMM/h/QOE1Ros+xwG/pXGCsMJW8BPRiTp3n
76XvwCHsX5VZCyljs9YiLIUrAWi49yUhUt4MzgJ/UNpWBMNdlOi0ud7j67kwSFyV0tCL9bJV/vSf
Fd+j/8jxuuw4SMHwrYP89NFJ6cN3aRiPJ/kd+17ovOSSCyFuFCzxT3q0RgtqPrvFAYaSqGzSM7je
H4F6i7reOOFdDCzccRPSFWb3wsi6uGhwWKd3Vu1tfvEOVPhnxwIm/JbYCyJhCMYRBlVnbx4KTd7J
4qcEk6e5qCVHLaph63vMip0H2PjG5ITotw1xpFHyHLFiXen7KcDgxN4qLNdfh8BXjaNgX2OhVyCH
MBZMHsF8Vt6Nc9wN+TviHd2Prb1dEFA1eD37L+IdNRufuleWuLJa8S16HcGDvdTXEw5cPF272AxT
P/osGEI4xqdT/Zem2h/41ThHq6gz8RT9ZcvWQnhjVoUFqngyBP3z3ZIsgRZfqLbvnHseem/rUrSM
biC4LP9QVNdG90fWm29M4SSsXCU/fNtmDmsqfn0qVg8vHu4sTCo+n9wVlbVtBtt2AbnRIM/N084a
WVGuxHeS3tdx1T35V/TQeURPfAy8U4z72MrySKRUPJV2qxvB6UnAQr/fptttaf1Ho7qEvPCdzMqy
hCDaL0SdO1MbAFw2eNpn0oQwMbNDNaeLMhN0ZMsrsuWaFJhVCN+j9A+D2rEengxsBGiB7486M1SM
19+7hqxl7GXzmiOwIilnYUDSQxnHt5SO9xvVUW/KwBeYtm6zG/XinD4MGWdt7GwO88QR2HrP5V3u
IZTtbGXW/rQb/rTMjCkrumcGJPdP9BeliYFifXTCb3BS5zukyPZ0dlvzznJ+0gOTyUUWG/Oro1kP
OGq2swO+S+2zxdInpZdEyrcG5PzfOkKsKenTqpfDU59KP1aZMEibyfTdzP7UpXan6qoe7cVXw7JR
bVH7d5Md7hrm+F6k7Z00oRNqQhOHzl0Bdlm6RUMwI8Q/94UT8OR5NCLVn1H7NQ++QBjdIw8fFFOE
VWNAYDqKQoMuEm5X5JYfQczzXZfZ0+9eszs+2oYFFjHGwlEXZQIv4XYI3Y+GSYdw6Hjsc+0+wDah
x3CAhcSCqVjILH+Y256Xa3pw1qoPFoeUBwNRIIeQ/y0ANaDPgYy62zLQ2lbm3UQDsTKAvdDiquTt
iqiZMJhrNG/GdkUgGTlRyi6EA7fThhJFwBTg0h02M9kKxqUG/s23LMwOPGWy+E3Jircnh4T4DWlF
KiajrJePtSYUKA1VPHZ80T/jhgnxGLlxIcbmhVosdybrTm2tqdsksFXdjUUiVY27tBGfLryEL7rc
OcHcpOZo3/IXke659ChsBmrahlNkmtDgf1uFJmxghmNJmZxXXcU1TDMhGA0qDZZOSksknpxwk8+A
LBGMciJgUwvwjxpHwJRtWBVUo7bXEbzPcDKK23I+WtNdRmVnWJLFydcSVIN062ziK9j2xmADJmr8
Z9LOscGy6nC1+SW82RTxd44IbIFf0hRM8vnhac2w9JEm3TmcD1fxc9Qr6eahRR1ZJi33V8bE6jKz
wqpYeuYdC4k4AclAlyGiGnMfiLr4x6mfDOocVnQjRjwUwQ0WcMzyhtDtlw4pUNtnrV0CbLd0Tbn1
wvBYT+EUlxjvjR7L03sZ1ujauPnbedZ7Yz5HwUjNVYCdbqM0zaXXBZp082AbcsptJV5drTbP8Cg8
byGfMAuj2U3cgIW5IUDkN7MRO6hqcnwWNfyoLCVQ+jvBlL0KdPILWTss1FSs5TBTJGgYvvtwetlZ
6zJTJJTkqLLmZ9PM6wiWv8DPCnri36Ts/PO4j2xSofY7cybWlqwXRdyCtGQ6DqJbJJcWDof0MIXv
brAAT7mtfe2EUyweaDWYDTj4ok/0kwTqFiCUGH0+03VBjtmItWTxCaIveDbv/JxbvCyAkRVmNAua
qryQZt/6eteds2OsrR0120aR9wO/rEVYDIGBMwZblV27zGQLTQb22Q31awS5JiWem/Nyai9ScHNQ
B3daa5gPW8vYpuaNXDptPEn3/N4JMB31xd61ODeTvvOTn45h5BkprjMhQ9B4Wk9D5kpkh/1v9wit
0xqSngPoGV1nQz4NHytXtq+4Y+8Wm3v6p3JuQ8C+T6LGf9FkidgfRY/3EwRVPG6NUN5L+8iam/yk
ZYTszUTpzsG4J0Y5SjWSqzvRveLrVq6w8G2O1NrRFzcP0QeWIGyTyYFxm6Dw3mYlapmuBDigezRP
KblAS+xHCDNuloGWbxXPjPhh5jrVRGPU6o89eLUM5q4seT0C5zoLQ6urv3B8tJETH7MVe7qEUL2E
eYqOIF8gvgZ8qEEBYFGQ79N3UjOtCaQC846mQPpop+pPLfkGG57rK0h7/eYPRm8hLpax4X1X60S6
/eqsc3sjTU1YD3jksBufza8N1JTpjnLFaD9XB6JLpLPRCpqKIMQ3PZdA4ijdr9rqs8x7lUHyJlJi
AG3baOSwEPtgGpvQUijVDxrUxeWcojsvQh3CBjxxou6O4hZ/CZNx8ns2R8/iC+1HQ1QrhyzojlcZ
Kya6hHkh6Qcj/++WvVAraf3hC606FBbxhg3+h58UFx5qLKEPxiIkWeTsPSV21BTLXmfFr+X7W9lu
lZnmM66BeM1UrxD9o7/k1/4Te2Y+z9ax7M53UYF+iYupmkq/onxRsSTnUv2jy1jFfBDAZNLfIEgF
HvtiJ79A3fdq6g9OW7Vgcb4PZpxQefUAwZ/UHc1obiEAaQ7D+jqtzkijI6e4SVdrVRKJ325Wql1n
s6xylYvb7qwAgXlCZDOEoMBhtLpBx0J5LxlGLeXp+TnwZFpQVUEP0ecsI315i9l0cheSBHC/+McI
9zUufDR1nRBSX9Ju33WABYETZd2Cu1jQI5kPNyQeOaaJRi0A8QnNaGaeRsjFBVGWjyInqoYengjd
th+Brjx/ytdDvbdS+ri9P3n0S9hCxyU2SvhqtXWep3rqY5bADbYLwzFAS+ojWIAoHpjfWPnfXTnO
WMui67P2ypJmbedlhsNV1anUMzbjyj9HYWYbnwat83kJOpulLG/Sbn3c52txCq+PEouBI0SRZSCv
Qz9We+XzjpJCxSmSjDHmgLMfXg+O4EGsG7dxH+ekailTQhPNOJEFP60hOinTFhzQhuiX1pNtzVxC
c7aN/TW74YTDgdzXANO92m561MPLqjfpTmuHQgwZ3tMlfYCvxnIOXdjTQaVn3I5OrSyvPGm3Wi3j
oGbdE1S/thTpbEEoXD0YyE/rYaMtkAq4DmIvEanqlhs6cAktnmUaQNZpAchR2UMKCsv7Vuj3/i29
+H3MgGd2jizCL2AQIaPvN8pVUBHOY9ts5yQNG+Y5mYZG7VDcB3DG/vm/ZkNPJ7IP71SlJ4QxxH1X
wkj4rCrPSZsuip7rwVPtOSmnR8jQKHq0x5jwVjJUgDET1iNHXUSbX5hh8b8kXFlx43FJJoWBcbon
IbHQ5h4hhKudOz3vSmFo7mKPyqztLplA7zvHX9vO3/y065VAjrtXplAz0iAWePGHYVr/4oFFPKtZ
kjCXV/9iX+240flybjnDchK6A6L8iTrG2nuxuOwr0UAGGrLC7jQS5ZSjQ30tEmAGysy5kFx8DeOL
AfcnuQdtH25iTwYDqO5lERztme/38gFWgV4CKGPNku/2HSeqnwsdtVl3tTCXmYw5UE9gaIN80Q4Q
CGWDf2URIoGCiaa8r7d0yUB0HSxRl+KTazmNlQ30ILM+GsfSytA787KOiQjYGdDG9VkJK/ZtVV9n
W8atqGraOm+8QxKfr/eu4G5y/9k7bwK7eqDvPKUE/Zn7/Mf1qyxQYpqY0HyjV88O2TVChVDJeI56
dZnsQc+nXYpSPTNYwc3WLZVvUgIPQZMuSSVmsRsSUr56GaRw9cc0qKPuG06uV+ndWnUDEmLLTsyD
uJN6Zbvk3PzkUR8Wl32aTUn2/Vt69abahdktPa5Je9TaoithQWjhYjQmZsk99wCWBEkIdvZ0PB4B
zSvLaNWtf/gcB2GT4VAOwt5mLc81d+FAmvh/NW4YVF0NPpaoh3zt6Ihot+rHvTkFQ05EaUJLVU2q
IzuWtOMyVy/agA6hDavaDzKLoF0YuYUlLV8U+XkYibFEzjVsIQTE17O8gxjxdy5cGb+9tZVvAYkI
zLJAymUyfRRMpVLfQwOCWF/9mvRv0N/MH3tAK9TeZFfGUJM0+XWZiNkvismNVNm1w0vyy9Uc6VgQ
JC05hvj/4QP0iXKQrIkIVn+yJyctV2RlSP5wKXe+Wkbg8n+9WJPnkIgX+nXFzsm9HHPQw4jQtpl6
I/wdTfhyYjrzQxUDTcJ2QVO8K9WYeq9CVd8oiWk5iDQPMR4QOVYLLhLal9ELQEnWhF3xR39vZxS5
Hw6RB1F2tp8orn1vSdvgnD4EXghFaw1lbBHurFUaLi5ErdUbDFaLWpQzByUoyAgz6JyhgmWl7Q76
/MwVp3teQnsvpJBtldPmv0PPL2AxvGgSVg6aYo/f07+6OUG7f5SdLl15F5S0c2TI2/H3LeIy2kES
7LUpQw86hjbUVsr+NjfOZDQKnehp52yykTvZyw1ZrIBT1v9cAg2rucbWBlK13NnTtaGSDGp6qWac
wf66Y2I7cbqqb8QbkCxxuv9K5K0fXfzYRYFcn5WB8s3sRchJFruu9Gy3hgk2FeS8fvQPsr4t+4vU
Sbqo3qYeeZc4rsJYumvDvnsPvHKrDaIHOzSJeYNY5DxrkoDkf1+zr4Un1/CbQ8FKBJhAGbVP8KzV
/o8rkeRpNjlldxUm+lUPTbFTFmk2+v21RcGyEnSBBAxKYgXO+GYCkHju74bmHk8tUgq5qIf6fxG5
/OQufIrmaFgIYZdYAhpA6a6yT4QfKB9XklCpSYqQW3anvLG7H/GPrbZI6m1wM4p3pw5zcbrnINhR
ZpPWZmfjacDlwnX8bZIP41XYBBqPcigBw6KIcmSfLieqpUmNlzJ1HCq9MNV1iiEchIngNbcZcjsE
Xy64GiB6kA/FcYWVW7djI/aYEYexy9x/ICVxVmVJHnTB37sv6TzAVqpaTJkWle5EhKDqMwqiaBHB
DyAWWm4YRZ0bezXNiWWAX8kRCrgmu/38H6jdaynt66GsnnUP7Dpjso59wfXYG6SiIL3MNe8fLEx4
Q8KMvEjeaWlreF44NASK5w1PRdWsq7INDceLK6b0/8j5S6R/dGAVyUzvGtkAwCFpxvJ1TYavwKpm
Ot+dr+OeOMRmfyRMugGru1q1lK7zc8i1xPhtU0uWd8usLASOC3+PSfrJCtjSx6UBmMMSS4/YC2L4
cCStzrI/GXtUMV8eF4zJa9wY6Nk4hS8tqKdHjGymMTdG8o9GJiXeVqfO+91YtiFLY3/iLa7CUpKW
iepPCKzoZS0Zr453kl3wanFtTQq17IaaN5EGegmxSRPbI6bOnssR9Bp+XXSElPGQAaKGyt2W0Z2y
DN1GiHo4LHEXfOFIqidUEYWznRrUofR542npzgE2ySLnLN6LqcRjIsUJ6Q3vJWN6pZIzKOkjZYN1
DX0Zt6NolgxHVw2gi14Loc/wzLcS/+kyXCFvig6S0Bf5cGzPxf302aQg7Ga8zV04Jg7E7NADp9r0
VcjcWtxeZYPMRrRoFEIohdZzsZ0vU9sVYSOURmSRb6NNUWzNb32bYHjZMglwee970QCWO+D1eHqh
viN2LdQUZkm2b86h4S5U1+mofsnAHo1MrayunVmtK/g3doTnPzOnfaU2glUAvgljI7OHES4z03D0
mZ9rCTE276je0XmnQc0MagNZ/JyfTRjAOcIfTnumGWrySzLGRZkT+vpA3tVzds4AOuW4ZXGhE4Z3
JpkQ/Yhh6OPI2qv3/y6zMaDEMpUk8FCtqBqDwtF4rUY0RgPr3VN3UHGrUmTmwnGdEtHV0sICk/IN
WQv91GY5jSsw4L0yk/kCgF5lsI09GHAHBV133tEh1iWyA9drQNegTR4/oovsDs4HQO79T0MixoGA
1uWNSEBBQeZjiPqH8O8aI5c0wmKHlpsPwal4z6DkFL1pBIio4AUYsBMDeynFeiOh6HEvfUbRM6W0
ZaACah2MkWRYg4YzyEU3dEOFhjpsDrOCZvAxS5p+kBGw5nMoh6grZLGTlE9tr2Zx+ypVMMyMrtu2
ui2yQ+7zQ6H8PCdfaqaZVh9VBM6GZIKHoQxvSo0msLShPLGUdY7gGA9OLVlODuIKg7WrbW1vtc8/
b/8bI2b5e0ok1KC+/Mevr78NmRrgZHuSKvqJGuWxsrhBT2cc6o0u4CFpmUtsmlc4GmDi3IhoMIaC
iB3cOdaBVshqlXBQJqH1Mfi6ZsFAnYBOagUKjFnVfdVelLj2QLs/CG7vK5KC59/WHnMD4V1zsajT
RVNBfiwlYMKwWwQ0WVqR1M7fC8Jw95S6Wv/DH/pUoEKNJkrEBo7wzUTovbpBJuUbya0Xvxb6otuX
6agFo/jdgkFPN9LH404nAObvlJ8HCQVunJ/2Kd9kYK/yG+Ng61mvorhgsiEpNdWhgQD3lVMOcxCv
KwqUqcLSHE08AZg1Ohsg4baryCZ5gFwr2SuW/8+lx5j8/qo1Ie3TaEZ37nqxQAm+KLgWBEu16DET
fIcdRqSpDwPnXXdJNkusr/KrDlOoqQTGeOopRf0wKTu+KW9rH9zcAjcw3viQluEAVbXXpskPxwDd
hYI8HoV8FsOOtTSMwpVHSIaHwxnI/j3QX4Yh+WTcVcYg9D/jgLGdzwCHg6JAzhR0lUgJPwJzJC4E
jlko/qm/hVloIHkc6FKRLqa4ALMPG8K4sdEUMdAWgWvmCFskRrYy+aSBsklPdbNOjujEz+Q6vBSd
ZTjiJ/8RvdED2l2T6uHs88uZ4BMboC1b7Mis7YHA+BGQLxosDrX3XQyPSlwIhGTt9+vYMpGMwExZ
YS7R1qV5s5pgXQXDhX8GNug9whrPMRyW06GKDZMTUFe/IO/PUzK2ihJv6o36S8gSb+0lChShyv3w
dcQx4lN2yaiJOdLnzcLtUDbdocKAERZTud9FFxWeRpgOzE696keZANiYqNeD8vmQ/2cIXIWnrJJf
wNi/wf6/UveLBXo5IWsAzmHviq/TLKyluygNZv3xemCk7RyZ8zV0qvR+L2aK8iVdsGvK7yybos1k
yoWjSeT4e7jiwtdJd0wcNI/wHGfVOo+7YYO6h7+bEUhzovunMt2wd7s/KFYX5jcemDNzArrafFs2
ivL1Kfh+PfzdU3Vo+PPIGWHv6LsfRmDCaWpB8gs39ywp4YeRh9YXAAg3UEFQFJSnG7hILnIK0R9k
8KEo/DlJFj7h0pEa0fWJlPXOAcwkTZNHPFKPEH/LWrQKt8imvaHJS9ldKFMUuHSQ/gMdbKjD4umx
HYfbdyFwL+i5AlmtKZE3U/xV0RZ02IZvtdn/bNjG7Ol1+fAhbzBSQGLZeqgPKQIWHOfnkmdQAIo0
wemt9JYm+LmbeafbSiSuF6bvRTHLnmlfpq2hOQENCqQXCme1500zcCoWjn6qf/z7vsAM+pfhCWQY
Bln2z+8OQYXny6XhHKM8+rG1B1pdDjfMPufuZMyu6YToDwMcXZS+ZgRtC8dbApZjD+mAuY4s8rBs
Y7KZ5reLiZt2HXcOhAxxikZSqMuLVTOgbW2MWtrqjG6J0k7iIGhD6lVAAGtL4PVBxtkI6E+UE6Kp
LnhxnnwbMJzEx8ndNIxuy8oDf/1NjlxCRev3zKdCpZJrSdoxsVlFCjsQESsUEXhCRudG6ntvaAMF
xmGD26Pv2RO65kJd+OmNd3HzDkbF8YZQbG8AQVFi8VZ6in7lOxGI2x0S9JKjqbLpLlCV/oHevRLL
EbB0Xy0nGkHQVHleendzbl00tFBrB0X3KbuvWbrThXgbdE1C9pZcK57osSf6myCkX+z3qx3PBEr/
USS2Ufbn9IEid9eManj5/KvyQt1ZBjCRd/8qMpmi1FWQm3oRy95wNnGmpnlNGdBLbMLx3mMnQ3FC
qnv7uwzO0sPLyypXKRC4sUtpjsaDfgZ+TFV8pmjYdCK/NzJ18eTvWvgFp2MC3EN7+wbUEY43zHkJ
ZrHO6C1Eik+bfc1HXvBMJW8TTwkrc4nnthIOxkIQCSMGzaGyDYA4D0k0Q/lqvlzMHYVqCMYl6OF4
iQL8/tj+a4z9no3xLBJhnOWCxfHZHg918Y4aZabC39cArnoIE1VI1nmt645UKc6iGSTIuoNseWny
7D7jfYiamFZZIWY+OK8xKvhYVdn733VoVia8BfVS5eU+s+JR5qZNv3kBgO3C6sZx5MtXRgbxqhvJ
Eugifocl+UpYHzARllXwO4W2H2cWFgfuibbhPQRf/g7aMd6ew7kdm+JU2oiF4D5up3pOvjhlwxPR
Dji1pwtfd+CT+stE7m0StFwe+o2s+Q8lo34R8xRTUSYKU/5bkLXG8EeH2rNhROjsWsAFqIUZZ6oW
sg6SKSLEMdczyUkOgytrvPN7ixqGReVf7NWeoyenf44HPYcTvJ8dKOZj1fMjx6RWnZf2vEXDRV+v
7Nv06x85+waTDv/hCL7uQpYfukBzDMxkjOLYXhB/5lWGWrR2TjtqQL91n2cCMWsAfOGcVKwZKwvE
IzokiFrZmrTVtoUH7BT46mmdwQdY77a9ddJnLL9XfAnPNQCLMbuEcLiXx8oUw7j1Hu8ZBhc4B53H
zlIas7QJ3rrEKw0iH1Y1BUC2rUOX9XX9+LQx5/5D26wArUgJ5DwjLl4LD+ZsohmgqB4WhlSGqbK5
FDDKPjaLitE2dmuCFtwQChTRun1dKM2av+eYjXufqG0hOuQ/YFrnwiMPuGvGIVOD7zNrcfc8tvt7
mVLckiN5yODU8Y4i/JsKmkaG3b3xDJ7VpuizHjK1ViXi0cIuJPxBqV2EK88g5HbpFSCmRZN4vI5x
SCdc/dmR/I4TcdN6Y+UeH8o8IxAaG2WppzJS4KH3mvfjjYdJ/8K1uemmSgwvHeMZhNZu4bGe/bU0
cHKS/U5WN/oaDxN+tlVTcwPUwvNLy2QpGjYCkRgWTMJ/T0fYzN0FjVU1h9kAg/JB24NJtSilLLBs
VIeZ2wE6LPCr03oCACxkEDpjEl88xfdS5SuIf0119RxBFUQelDvzV1rBz2tbq9bvRfp2g6ltkT3p
UNtlzMb9plWI86WlYeLG2BAUKBgZPu6pQ9fxaAlU/YY7jSaKQpk/XC56B/yvXCItx+6UqDN4e2B2
Alg7OFYeDvtrKtei1fW3fQ7l6bgmLQGlreHyennpdUtoGoPh6euhY3515kSy4eD2TC4CoRy/ePUt
e7SRWYIwALyhHjqIG25hW77cPS6Fyvczx3Vkmj+X6lnC2vQT5SX+On8L5aSww5kQpWYEs0f0Gtlo
VLUd7IH4+6sl6Lijm16/scWZGWgedVc/bVKJHHl5o7/U7tLr59+PCOlVp0kCOwnxtVlQ8s1YHfBM
uFm0cVvxF8uDrz2Dymoohb2PuZEF1Li2HlbkEbj35gx2L91BGzRIKYXXaP+dp2QdslLuIaD7bKWE
irt/vhKpyc2SmTZbuK2kIRuHY/RggfX4UNI78aHyyq34lcdlKCMIn4AWy7OhU/PXRci2lOS2gidT
l4z8/caI140ksihhVWWDrQKaau4VEWwx5LAdzPr5xCe3sJF8IAWdPYlEuNLeNyIidVJuHPlaP3Ez
/tEWc77SUidl7NCaCNnMWjpw9874RGms8+Xs9XcqQQkHz1B1rJpnc9iQlAhRUESI9xLnhmz2tfsv
7lMIeGAobZ6pwNFs1ThwkHQVKr4aaZDJIM0vG0IXfThm68aKojw7yAiXDng3ioCwrAH8AozXRruf
jEqCKebHYU2cNEYLGIxLYLPTGHuWy/lIrovac3mzFH5lMj2aedwwBCeP1grS31KQRIwTI1Y7kqq4
tmPP9ljzWnCAlVQ4hVtc3ipKtm37PmdQ9QN9U8n7kJBPXOKTLUsA2VatvJqAr+G6xvTlTgENbxnY
B4hZ4L1+nz+oiod7kXnrInAJOoLbcsyoiXsdRbrFIWRXLwSBLg68DfHjn2rBJWJQ9SCTOcwB5gkq
vy1HEXoi71/q+5ioXPquoaCRF+ivROPrP5WgxyInuv96+4dTC5x8ifS1zZhwO0JWuganSqyHhjL9
XSsOhUSoeB+gFJQsWNJt+9EQ7MccKvXbQBEUgnGK1DRruRCzEwTvTlU0MwNzzUH3EUrrFvnY7Tu9
jtuHIy7R/yOV24DO9LkMjt1nUqyGvE7Iv7ucGhPyig5nj+9WP1mLa83ivQix8f07iZ6BDD55A+8x
BvwQcspbBwo9+kaBHt8mQZFV3XbDNlf5COkJ/9QJnJh9PBRz2uv1jbFoPsTgAG6X5N/kb4+FKjoi
GWbuxIwTYzBUERC+Bw8G4dwb0vUyqN23t4JNO/G9HUVntuZaQJHc2pohKp7UzoKTlT4xzyXOul2Z
xKs6aroUlbCz+9JeA+mPopw7uKpfkOIsTzLZ/UowAcsiZ0GrkhmXnhFz8Mt0yL4P/6FteeXErwVl
Rvqc0CZFg8BrZegKuVijVHxEetHyDBzccq39FXrvtk4Dj6080qGMLICXmDg4TKJOQZlJUelbGwq+
2+iN9yM73r0ER1XfIZDvlfaCpJv+XYqYHiH+w9m13VUSg1hTQ5+YlzCgpDqSFe1SslWCQeX6IHbz
ASJr9aOnCbJ+8j3io9+DJa6sxIvqqIOFkNlRGJj/HTVVXi9MquOL7vlq1b0i6IPSygS05xLt1/i6
Tn1V6i+5JiVwyv9e2KALsPID9FVUQ+GcfiDTg5dm6IxHRnIY+W5idiOVvuTHEL7U4DNfoiPdJKEm
ci3iKW+U0iwNpZJ9Jm1HLVjka2lk4giBSYymVvv7UP1hvQWmuqWB/QzoxldBv0nlXcoxnCZz0CDI
UsmmY8ydIYrpVWA9USu6PXUYDgtZDfLBh8HPUBYgQCuSFla2QPxGNi22+OIAiFA6lmYXDx7I6oXo
LpjfPBxFjMUigBfbmCI2R1hJzvX7p2Wbh6If52ymutho709t0y5AVczMw9Z6T9DSYw2p/LqK+Q0x
hGaGi7nvXbGzc6AbbyEU8mfYeNHwD/aSpA4iob6Lr+muEn2hywu63BPUFqXqkWt+joMHzXAO3RrK
fHRG6XbKqg58K/lNcvvkYSWuTnQbyooP/+Ryuss7WNZmj3Lb+xBT0PSZc4upIP9US9udRSKfx1ym
PP5TeQgSaJa7YPDbjLOSXMlNPNf3fta4T6kYoo40PVmYK/isFsadW9CieG3/JVsaRTTAgnMcs+m2
ACRybjDHYi05SIEm4PoXzwJa9bMGS1Lz5SXO6VUBLoMrDhCdmSVBKMt+wbPtoYFug0n7R4POHObO
M2jIdc95AVsfkvZXRxAQmWqJy1XxqYdNfujjBXIyrtuKEMFJRVF93RDXzWIqTTv++79P8MRBkxPr
0v9Q67k8FaarxRgWir2qLLyNDSaP3MpghOO0Uc7LaHf97M1gHLmR8K8EB1moLF85k7vtVUUFGdUe
tzDoph6Tns4DQEsem0xwkYanv2D2OsaP01VXcJMWQeget+HvRipkCuw1NRTycA/PKXitFMq2cDtO
wft67JIsEO4tvBud+bdO9qg8V7n2fH3wJkVCKh/LqcGJIfUwuMpugejSKAIJcwZR/9syTiI+D3cu
PTW637pfctovNzUjvsc3dLSi10BJHbrK1C0z/XHMGZZW4OE2jMCYsh4ufPhUdqLEhMNylfcVXa7e
+zN9VLH86+8N27yvdcftM13LjHy5KMX0I4QHMDKSMhp3YE+0uUKHgS2UFnbWx+uAlRc1CkRv1sM2
eqYMYmDWFaOEjrzV8h5AFFdcepps2D4HSAWhRKKX8MtuKAlqm9kkQq24V/EY5kihM862K0Ohb3NU
WCbG22WOqDgsq11Squl38hcvI/pJNVYMJvS4e9CkTdAje+dTeXtHy6K4oY9hgyyb5GWlUowijhCv
bheV5z1EaLZo315qeH/6gHFNkhcIlRNzsOtlCXMItY/da7n/35zixa28Fjz4LX7ygjC6aMd2yPC1
Y0T/wksg5HYmrsEZ/EuGrnFyuFnsjTZa2beoqwXcBrQADerDHHgSQ+bJYIIoAIzqQs3C60QO/brN
0fCDCysZ0phS/WH3eL+gBddNIDi4k1Det97jzz10/RkxkRwiVY5vDurTGSMbb6MUSG1MrdMDozvk
bch88DjVUUqJEd6aABgcHp58w2umrUurRyWR0/n8uqvgxAwLFAKhXQ/r2dgACIi/F7JjZH7wTt7h
I1xA63pf1p9wVy8DLT/oM5cXpNgLzO7rRc0pYVIEKlNdzXNwD/QG5BAxTTo6zr8w9gjELudv/A//
gdQ+1kZBlREAGrdvgMePE94Doc2sd/6PLE07EHUnGcQM8cw3EgBqpqEdM9LEs5huWJrAb5/ScdlV
rYE7WtMT0vcSCD8neEGeAD9euVxNMsYjaI0F5tvxGPIf6P+8wyvHiCsN9iQJeJZiI5y1lDVDqgJ9
OY2Xa8lj8/9XdKU5k/MlyqlA5GKA1pcH4JBxDSf87CJu0VdidEqjarhyYQlLwVHAmERVsVlYsFBe
Kz2dYnkdRxvL/+Dm1iPvwnsGm4z0oJ7uEf6Dh59XL37CkcE/13u2S3EV+qaTMfF5GV41hRn7+pl6
WTDvKwIgh4V68ad4lQDlhRnAfID92HIJddHNG/hZIN7bhj+lK5CKedi8qZt/r65t3L9EkAHcHeZb
aClOpV+/ln2qJXpakC689ympGY+hPBP30T/Z88OradQ5PXo0aFYDtjnui31Ch6GwPeZeisXktN2N
ZUU8mVMoBl0dybOWKG3BtBzN0f8mW+VIvDxKmeHxzVc2S76YPC1dm6JdjGpQIcb1u/re8080Chfw
J8wP7OPWxQ+zipjr9h7D/fGjEeoBqECnw211AMH+gJoLdFD112qVx8hiZxMSTmh6NAXgzrqKkwhv
r+9j0FGBYSo/o2uYtjCWJ8OYWkppq06UBVu5DQmUIEyRUyGNdCCuS+07rpkpbZxHdcY34WIhwiKe
9EhB+9vitrSosZ8oEtzs3AR49zPhpo49VrN1trgnCrWfs20FZyIkHkMBvcLEQSmKRrR68j+Gtayl
R6u6CKPH95IYXOovF+mqPjh+UHwUG+NAVc9OtQ++URUVacC9nOBTw0fy99U62yBhsGkm7+S2P7+q
btMgnrxli2hbjsXLZa4P4nV9bNQUlL43sAbR+z+PY2Yu4129RmFUIBeNaSFpQoGNpVbsBEEljjjy
alPnSAdvZhDMyuDGGHkWIoSlUEoNlhGOLEbVqZcLIJJ1J3rt4JMd06EMArfdvLP5zaaNj4xcWUZd
hCnmB+OqdBSyi+tjFMPo7Iqu9DFWlN/PAtUcZlGLvIJQWtA2c6upDdadced0H5XbzxBZi3hoVmR4
5Z+A5IabuPW490AfeX9M8UBr06n3p5ovUTUfob/SI8t17tKnLU4wziVrYMUlvVciRsI7jNN1Ri6S
chYhkkrRI9ON88No1SZsU+7maoTOqeYI5FMtk3W8moW4x9uCl7HstXJYCcZ0Nk6UjkilTf+MM595
N/JmQ/pAu6JUVzZaDtgv74hZDRk3UugO4sGsD5bilIBngrT31CO7MGnW14mVH1RIT4YGtxImpfpC
q8BLu+UfK3DPc10p6pLnB6/u5deljqakiov6ZujNbk9spl7O+tVB1CdmV0H8MylFrLYnF7m6w8WX
0IJwZrBrd7ootG5pgP2HsBt0QxUTrZwyZQgBEBQ4Vs8GDkpzqif0NRwNv2ULxeTVhF8RAiXVIDoz
Ocld1qTmybVGp9oqC91Z/bdmMgv/dnXdgyoUPcuZ2U1Vzjg622nkj/6ZEUsdjbbmnMTnp1q0jGAE
zf5+qThMWr7SuxqqSlWWKOar1iv6TbqmJ2H7g3y6LBTCfSOje+QfHGvqahZfbpDvr6FuuoMgXxUW
m3CAZC3ZAZovIxkoWTS57m2J/pydgnWx/CQk5RYRYtERHkcZGo1y1iagN8MPtBP99S9K+skV9/0D
SilsRX5hBDYvSbMTrmpY8RTCtFb9qd0tBZoAyn9SflY94X0y6d4AJDjjTivOCMJTjw7Jp1ZP86gx
YLLzCiYwsbwthecMnMCyLYJ5OpUVPgy0J4ZX3rQn4suYkpn6GyLpk9syn9lX5dNtXqJ8uPOHwOPW
VoMiipmv/ffE36sVZePu6P4DqdQEIapf+Fw3ecbNkFMR6MbNZdGMaOUUqs82eytZ+XTjVkuV5OQZ
Pmt9MTWpwxOTnqoqlOVPYUt/5Hb0KGLIsPboCojNS1OniG/OsedPjpVKEZjVrERWpBJ8HEmaG1r1
obA9w4r89IrKK+0bwNVTmgTcLWN8elde7gbHrX32PwpPhfXivmYbrThyXFP2X4dI2xy+WATZgs6g
cV43HXAxDYvIpEQEbgHo87uffj19qbIMnlB8BVS4vZwd4Rt1o/qg82CXuBJdYBJYv4IWbnMybmwS
ZWKnr66k7IEi1hrudCu7p9S5zHgKunrxwbXvcsFd8mLw33VqBiCy4uUB3GgqznHtV3Qp92AzuaKl
5EbNI/nI4p9ySe9IpUd1GIdK70/hOAzQuugvvPnpT2UXhQlFijjbol2QvxRKfqnR1WoZcdGcX+Ma
JtYyJsxbJ6tKoX8iQgsa3mYl+UZ9g4R19DMJdgo3cw8hNJI780ynJkJeV+2fCdtDg1zC54UPxAlN
+Gb3VDP6uMHaiP3WeFZy6MtRb6WwB1f0Z7yr8mPWywE0ic7jKLLcI6ad2OI2ErZ5mvrzRKhzSlc1
yJW6lmf7Thm6DVjsN+WQN9IIM4fRtXwqH8B+5kK8WyFQPEPgxL4jpyV206y7j9a6ZEFA8tvppIKj
J/6HpoR+EtbXkmb2epoeKjEM35si6pOjQpPN1cLz36Z5k5T6BgPdhnrA5xIQrPyzys/yAK6s1g8z
dFcy9Z3WPE+4baeZCxylzisRddvbqgPYaAgQ2Aa5UruvxW0VsnUIJM1xrlQ+QNEsR9ewwKEgLUI5
VLjH8IZknkOLJoZfuT0gIK9QdM3MyeGTZi/h7Q+LOtlWxZ2lrVJaVQgjxbSX1YHz/88ouwIz1Lnv
gu2Z0k8cPz9sa3kJJIUTzGVbNqmT0vGXCFfLzJ65SiQTszaddDjwjz6V2RF6wn1uG/7FogeSj/ye
fS89w0KZWgjP/H0/RiEONSiTxB9CDchcgcVlesYVXqrqiJWsaRW8PlSbS59M5cxYGezbf/NNDDk5
lnMpirGR1Gnr8tXmSnrk/mcS4Bi7fBUrhJQN6az6oAHPC25GIkS6cEvsEXOOnYju3EsImPu7/rBP
IHJmcZ0/Cl2ITZ2wy/uhjZwYJVP156rAyQ8jROfaV6XBUwHxj40bwcJ3XzmqF9+TZbIBL6W1KW89
CiWYjHtvMZd4x/op0bx/WWX7FRtyX6XQI5aCUli7Y8/CWG69S9bgD/yy0EUKPvTrX5dXlT/uXWyg
61toye5d4ADihcdrzh14WS/WWfXlmGOiLQBooe7p8XdFHpQfxw3pOPKKEaH3LS4Ko/WFB6rfz3UH
QtxbfnVQuyqWXOwkhIyzD13ZibmtTjCG1WcI4yYYAEsrIWDC5MYcKlacLG4gZtttGTwriFFcQTUz
MopbpLw2Ipwmd5AhwCmo3ppblOtrJzONspARudVzZd+2tLySkeXaHrepLB/2uNg2gpmIZyyYm8gR
rx8ux1rlM3ST/WnSERj36hy6x2Ml/LJcIj8/267RBRsT7gyvERzzB8b9cRRCTDoN4N/0SrC7nmSk
3ZP9lnhsTi5ld5U7keFxSdqDMgF2+WgL4ZMky++U+nT0cWOWt3ktAJUV/usKBWtZab9PId4ZZjVr
ItMVQOOlk/l7N7yLT9tO3vRH+pEauADGAEwIg6HUn2/SU/eCG8ePsEKYxhcsS6RAWQZEeAIoM8RH
mOs0BgAtJ/yhj/+rX7Og3ClYl7cieVFmktOiS4KLm1HcUxT3pLKeKA2+VL3DQ3bWDJfacCjVBrT3
DKgg9TyB4i85pqp+rdIj04c6nC/ndbuATlr9yU3ra/LyztcvPKghnAXvEUostIAHk7SRB2HkPA4C
wZJ/AQRYwgjegS7FaxsmkzUM9CFa8eRDAwhMYQKbhF38FNvDxGqJeaG/0bjLXuDauOprO8v96ZCU
R9uidaMYJQaM5riVP3U9goyj8s9UxV6Syg+N82NtaMLAGmylPPq871ovK3IoxFlfz9x66Ih3fxkt
3jiKb4QCs1H9da0yq4odo1DRdbAOpeg7M+87WmcrfUqXY5gQRcZYqQJwsWOxw2b/CeBEz0CaKLXQ
LlB0H3GxEi51Fr4VU6cdMUjRO1v0Ilcg8agP1bvv0UWEN1/kcxY9GpTzGL47Ug94eApP6A8/HCfd
dty5RhYM8SltNyNcsULK9GBpgydp0fiHOUZ4XmaZkWxg7stGuUIV4ADdPmHWv8UaYRTQG3wvPDlU
KLaCAIG8w7qz3BL8mydvi/5x/UMBsGkvI7uXPWLsIdWiQMppz2ZXCrBnsNlC8jEK8wi1+C0LRjw9
TPEIUJ8vQI0v9gZvkMuO7qExv/Y++oe3FXn3LzMnSo9HGogt9WQViiFSfItw9BwpguS3/rgb9N4g
TeCMf6H43PFa4BtLtHbp5d20x/L1TGRHvwYfcAOVnqaZ5aajjaLEkbS0z5CxIHe++ro7oKtDgjk0
x7fGNAqd9YHVGQna+zRhPEJL1yHT8iXnzQcX3qwaVrxEN/tWYU2M86oxRZIPZaC9vfv3OJkYHgBg
cimG/PSnoUHbPS1YiHwXvEUu1m/jx6wY/oOKzmK/RErkeZAhdjSfJKx1ZfYN3CzfI4tb0KiEEXGI
NuqVNatE6p0dY+fMqHgQ4gva+3xYwxXyaU4ksiuLDdlwtMatjOJ4Ks5KZISE/XUCR2OHa52Idfpv
TsQ4mK3Js5IHLVUD5TjkHCsxyoCeAGjihPTj7g9pp9oC2pvTXirpOkzV/JlEnYpTWsy5tHhaeoXx
R6RekwaCv7+RrzZJ2/m0RFy8LxiHK4MEDTo2K9nL4mn8rW/IXPOvLR4Lq8xhzOzr35WEgONBmUKM
nbk45SbCElWKIwxWUS+OTvhu1gPclSgg61tsCZim3ubmfKgFv2EPGOqDcs9YPOvlDB4aG4ADIPdL
CXxlriciiuDN8XgS5AQMyJVs377eQmluln0THj1ZNtCvFCOCkrCW3QyV7EiO9bOhcWM76AHvNbkr
uDihSnn6eoYj4kyoP7G1IAfIRqBiAabLZV9wZrY/y/yLd4UzH1Opm8/lIwxe2wrMFZ0NU2iVRGIq
Ix4uOdJ6Z6ajyzF+IjrGvPr+fNuyj5jT6+GHqVvjUOKhkEy+Ic79ewDotL2n80nRubIDXX6tv6+F
IAhf9Yifypm1kXBTdOscRcd80gj1XuiXZ9SdKplCLf4oMAUV8Sfi9c3KwhBNshTzbXgOCzYVkwLc
D0qdG9soqSUfHNQUZj5YrsqXEpdb/0usIJF0qTZn5zi2qR3DdkheHsrZsjkgXZ65q0wNsGel30sU
i1eQgTXORKEQrcymLUMAshYZgligd7OJBsD1Tl7tUYq/V0rJKEp0ixp9Ryq7GTwa7jNTBYy9eBTI
dUptKt6h8B8zjc6QjCqu0IANlJ+sOzw2T9wNNp8U5DXhUDlEGOjDR85wblRc4a+UrmgtuQzKFxYn
zO0QURerGUu116j1a67tEU19KUz6u4rjLf4HMQcRgjKiPTdRnEuADX+XGNQSOmP4a7ELyF2YDQ2e
KS2Fi4TRQ/KNlc+VtRD8bYlhxXMIcKgBWxJc+ioY2P2rRBJRkR/LDmwMaQgOCAGfO8zHv0OGx53l
32/pzyGrlwz0UAn+9or22vVtDA3cqVbyXf8iIecKDAIZ+A1S1SQCJ5OAJLEtl+wpc5/RH9eG+JKT
MENXdmQVooWaRLA/vEV0eSWRezAjkpK7047A08Ek3Z2jLNm9jftywWkLSn1Xs5N8Nr54MDRJk7qE
M32597M66rKdqHLCAcV2zQvsr2+pmnHOfa/gz0Mshr1a453VBTKeY6sPrUo2TXSuW5NY9YoJJ0ke
R28nTkpkQMCqaXk/FcO7uSrvXeBUanhSUGjdmP+8n1i/XZkhP0WtlzWNjrNL6B6naW4N3XZxiUk1
h8vd2Eo+sTKgVa3x4FW2xfHVRUt+4V0AWyBf0GkInDwnEA/POyKfwyJ6/zjc81CJqBXfvfo9xdc9
r+Zrq9a3xquMDWpPtM21bfXLs31sMe20wWDSV4EjbJFCkAheqz0k1/Z3f3XOdu7WLyfAs0Vheg/M
DOU8H6tprkc680K1K+lEL1ur0q3mN1DOaGAfOpuym1mp70Bz+ho/3hXfLjtXx4593rISl9h7K4i3
mq7D4SFDXe6PiyauVJkehZkSxX/GNsv4pTgnPa2zhLo/22ZkPd4t3hqDxXPCogGr9UP0zKti8HAe
EzoIoSqogSr8/yZ/mC/t1JTFzxJiFcUkuWlA+dbWiKIziYepl2BkPrB8OsK5QLxHbguhMU6wvAEq
+KyF8v3trpdBq2gv0ssZa4UIt44fJ26F9pPLmP82EJZ/vA3SPNcLxSBHzfSYat6kRaENFG3uM61E
HwmBJt/BzE4Uvch44vw6VuMJqKbTGS1HXGUg2XVSXuHRzlOxTk0sTdPfYOsFiHzTEJgaPo3aYFps
Zjy0UX02LeOWHkPbL22NEbggE8wDfMO0efAXEOKi0ZsA10nHNg+/SC3G+dfklV7L747sM6DdSQNH
zYoYkHXGwZRSIKNscUmkfr3FfOvp2KcXDQBs+9e+3BA/a9iGWoFP6s7mKgq6tMNS4YtCz8f7aQ+N
DtyUdAW4L708dbIDG9PLhvJTy434rcUbOPvUxauOren0YwV09vvF/ILfhUvj3HVQTya6tcwDdErF
zopzOkLZjDe+2hJVQO9ellNnpWtiSlf2mnJ9OGGykFTOVs3Hh+yAt4uSSu9SpzYaafAjcjfklKLS
0cAqgAw8uQ847S3egu0Xrx4Itt2FXK876aAmm4op8bWR8mf0JEXCx7Yxwgjsj4Ekh+grALtE1Z9Z
bJTZYbA0JP6Tx3EU7REtqUAFfOW8y0HCjSv2hRux53rWE/AGgV3UJwZgvQvxfFxcn/wByDSHfaID
2SAzDtW7MD5Jimc/4zvBZ1mJstuum0TU1e6g/4cT/nZJKluEUasGT9TwF7qbTZqknczvSfEhEB25
b8y6qEwrRHhvZLlVwL17aMDMlx8Hd47/qP3TQfmRVRME3TTXVKgKKDxgztGQ05HnQm9kn4dH9fT8
pF5hhVIXspI7GtL4+x3hW+crcLs1lcSAsau/lDcdw7ULkKecAcSJV9CbRN7q6rVqomykw/q8Tmjk
iubxxuG9MBkM45DDkbzjiClvR6vuYcBpkKifVo3Fazf4a9RCLkZhf+3k2ZoBAAtO6jIISG6v0vcP
NO7vtagyu0GuBJEjeGEa9vl9Pr3RAkGEzLni/D/PHycHjPQnrCqBycZiTjpgH04FEVt9deh69WeW
cN2YZq9IR077V2EU26n+58N9ssczQHopvRNX2P1zmkqkr6ctx1mjMt04f0J51FrZ6DBsGqfJtVCb
kwpALaPp3wXlVY+JXXmF2KrKohlTEl3IdxgK6vVbWvi/P5vreiFzPzicywA7or/QrpsPYcX2XUOj
QBpwlfmysmSwBz03u4zryzDu5CPYy8soz6laYt5+6W1doEgyW36cJRZwFW9SwzR31Vvp/2Hthy91
0g7GtpT4U0GAIpN78dEjGKHvz0JtQStLdqJ2JUXG0ozV0CgTaE1E0xEtZvy7VW2qZssW73vzffmi
un2IjBJbmbPmP7w48quZR3yMWju0Aqo1CcTb5RfweeSit+mKWG7NiXpZRascrjPvcwbxxLDB/xPM
1fxLK9UxiWKsq2GQM4yFOp4TV1t+bp1QhMJFAA7so6hWW95HGF5lmt4YFemYjjSZ4GqeVKToNdrP
ZPIk/sfO+NWRY24vAwu3f3gCEfgBHJjZ934TCreOddKJ86PzZuJo/F9M1yH57d5+ReH2zCPtov8D
jn9OPFEnf0WEw8l8/6JTy44PEdoVldVXzxCTvUkQlbeau9czVT6nNmXSyHDnGtSEEZ8dHaNTj7pp
OXRxrWTTVWVLt8fNVkVSDFNXU54HtYNKv87n5cfb/rAF5ujpUHYcuGdBWCDn4Ao4/jljK1ttyfgy
/2xgfCCHNfC4eMTJmbkEQGE9IxoZMt+U1KdInNz4SBOzvAgCg9Csxfm7GOSQMNc4Nq+wFQMNAgJd
zWZb19pXOqZezsyYpx/8hocKqzE1r44wCLMJyQbBslGR2jmdCJ7swULjk88OB4PjkFnD6lW0teyG
7cNUA+11NoRY0BTHGtqtKQZkOkGBz4LcVsKhRYODe5cyKYNC8hCW/sHDGZCevl/UUNpsKBRk6HKc
dOO31NCIa14gM9pD5btP8poRseZEML729XSJLZRD3GxFu7AaomkW/yBZSFtPsCD4AttGVpQeYtud
VocM/8Prl7GKh8RF9nrY06lf+zkSqbmtJVZBdyW7IkxkNHBvZOlc9nDV2anFXA0rrQNQCwyTmwsF
KNcdtijuqq6AnF4BPann893Ulc6llOfpbuQG+KnV/BWK/A/fHEqxEBV/Z3gV/UIxdJWUwjGst/4U
7va3RnNrEq4wmgt0ztDuFqRxiaU74zwBqzy9jeilXGcJHjjF4Afu40MQVNmjbC0Z/TjbaGB5eN4z
gHn63m1qSfhKNAkp919uUlXQcwTBsxPBDYgdSeKRtcszye6pLhbaYHYN235g7GwWnFHMxAteUJ16
Y+lMgJtn6bQvFXoie7F7r+Dt6ubFU+3q1XF+UrxLdr7mWhWpMi2ft8FQyPQwenbO4TUxs8kPoBzQ
AxJVcbALjll2pvZ5Yjh6BAxlZMH4jrCmrX36vTQ+/EF3WPaJf6umRWz96HqQqAtDIyNYs2WGrR8l
aMjHDkcKZWGKvj8bl9E/bjuTJAd2+9b/hEcjDdhrvTqcEasSixEJVMNuK3lA5jJOwB/5Z0fNzTHW
sEI+9dtuuDVTA2oZiBtNwYRqLr33dZ0FnjOsSEpDYlYIYdhaSph67RuL4gLoUHkedheS0o0yOWDQ
ya31piM6122jIeBKjlI+vuCbbMgGvPWJGPMmYqh7deu7DJsmSYUkYlzlnqzJzByIOAJ1BrLr33Bc
EAKDZ3mN2C7Ea/u1KBKNTg1X1ODRniAqUdulENnGu60iMket27BMlQmYg26JhkG4zvU5B1BXP9qb
AtkpNYArT4U4CSCWs0p7Wjb4UO4fGDJkAaTSr0zs9HKhhwS3OMDZTs6EKpvqSsb6HtJxLv4Tf25N
r6Ll06lXgFS8afRIfuG0A2ltxPdkNKNw3rNDGE14N5YjO81kjBuSi6DRZTFgTOtMFC6J+/aM/0xk
DHfSLB5JPwnrg/Veb6fBSZsVSnqgxZMwmhczvOuOs0QSs5SWJyono/X2UaPg4ovehI1uQPth7lN/
UFpN2iUmWzHTH649aNW6vc92Z+pqF9cNbksGVwNpQTF4Tm9tJeBto5WQwB/7FeOfplAgolDEK+qP
UALrk/LlJ4qAMEpotoh75DzfdJUigkDeORHTTDN8yQSjnE1APmxzwjP+ZPLu9wmpsjOeXa0ir26M
NoDFKohCP9f213LWt3EjYIOP5XyBUXKu1sMjzhHg/aQf7Ivv3TAZAABmso+luQ3XHaoWpmY3H6YK
yMf1GtQA3tO3c1E6OJxZkoHPUJU8PTVyR4ISNNj7riIreYeT0AVtr3eRzvEynGqyEJZn4c7G4GCL
lqKzuRxMrgsk4QlqMv6xXg0gJL4Fh4TRfIMa5wPwvH7c/3RC4krBrnCgH9KNu9nuZgB+VDd5vxgg
bjZaqMbWrA7IOpzn5S1+a2MvKmnMT8mTqsVCiClOpllCgh0sdZ+6QTf6n58GsTs/4t4KnX757n4x
DCbfIqQMiazvehSBQfFegKhhP61P8PEN+slGwBi65vsZkVNpj+vBWK9RPYAUOyB6Y3LTTDqkOYCf
rCH86ubg6X7vSDiJk1rjIN9EvLlLQ/OoKQNWDrICl/6byM7Ki359ge16+HY+f9MkuvOTEu962Ls9
SaN40/q5YiYeMYrnc8EMZ7JJw24zIBpe9/5xgM0hD07bjW5xlJys0nNaIDfrQ/DD/QkDVxEXh5j+
mYqO3Efa2ChY1bSdQT5iR3pGJwsODLuF7c2FtGymHDo/7xuyedYGsthZTUGfTW42G69r/95EOj6A
R5InzPc5qazasEbShUAGc7B0N7GevWuiQ0l06ulpdjWuehcQgZbmXwzSSyATvx/+uUQgRc0nWRO0
YtUND57uBGORsDGUorCSJk73Oro3dnLfUjsQv9ebJBgoNh3fJk9nT6cURr9lztjfiwVhJMhjRRsA
21mchSwIf9iPcDpAYKfXlBc/RTfI/8T54HwM9my5cLHYWuhJPZffN3jhHQKakA4IjirXK3H65F+X
E0pRbzpvdPNgq2niFRdYtWqxyscTHKb6HPpE9FrqWXHGLJSGXmCZI71LTDVgoiEcPN9hZl66cJRV
YdhVL/6S7awMyz+p0nIXq6xY9DtY31KueK4M0pKxa/bBzcy71Zky9MLoeCpzf5etyrKt+YAPRSFR
ZyGUtX+dKjZV1Pl2XbRafcU2koK3IQu/lGBOiVMOJg9rYwW9qfkRddRnPVR1j26fnz0kJDaWqu9M
fJnIX20Kw4Sn5gWRePZsJ9LsUDebSsOQ9xxnDm0nyfsKUr/I/tOU9LQRoJbWtACgromEx7ghYQvR
MbQvJyN01IfIf+sLgxWZ5/3oHHJ3B6qmM7sBzycdgmUKH/sANkNLeJTn+Rf2/SNmcyxBrj6iIZON
XYAxjcC3jfw9Jt+Pz2Q+F2cCl9lQxrTvaRvO5WIyyQy/KUQM4XDixunXTOYOm2GvKx11URykDmRP
4CGO+DpB6VhNTrPgAeA1rpbzXRX/MuMRmG9wy2sfuRJL+mTeIUJpnHvy0xyYYznwWcPdE3vdEzzW
LfQ+N5IqsoCja73yqbFJ9nKH+ged5+J2Y5uzn9Tv2dGoOYTOZe5+Ei060Z//toqd1wQCN1Ld2izS
PBJKWeNekb7lAAunf0/0fB3t283nxAQ8E/CC42KGXxABt+2NHB9R11qHWkdZVqma4WlG+G7PIJ9T
8YAU9/JScmDgZ/6dukWjeMBSTsGch+ZFCidNrwM+ob+LD7veivrKbn4e6Hd8H0I9ky/zmMlTaxp1
Uz59mWsB3XNFANaZDGwss63wveDr4TG8F4MDZwKpiBJ1N4WK/jss6YzH1+6PzXwc5q86tEsZraxX
PRZigDRcaV0t0vlUNyOnwMOlQd8r10oXs79IchAEQb9aYHyvdh20+fK0IzAkyzQO3rLNOl1s7U+s
NUzgkfSto8Nq4KKxnUyRHlUPY0XwtM4Cs4AyRnbVhQ6ZskxgZ6PfUS3tZjrvR9ZYP/86H+HXQ7zO
Xrwij2I9EhlTPX2D2FY01scrRk+sHxXqOK0Tb4jZsvqRjBeuKnbrFlVkqJBkNYeqeNKpx+66ytJa
HiLah5/a1SG9n289rWyN8ygCHbJyt88YksJia05b90Fm5XIb4benEsMDFRdy/vasUu3hw6aQoJhd
cXoiFZuN/zlAt2nVAsXiw54pwP91idcmKBniZIcfdJ0Fc8uHnTk60kQkfP7OIQcxA5ekS6kNz6QB
8Pp6qllNuWefagMf5H/U/zi3vVFvumS2b5wx02+G8cYPsu6tFsi/AWivGT02F06ILkI2GUyh6cAh
g71BAJsP+Q90U1iwZTzjD2WETw/nrjoUAJw03R8G+LFWUHzsBYUKx4KKLoUpSTMVW97T2LrZJ80x
+r8PbS7pdvBO42VrKEIdHdPrzgnMtzqsI0NJlgiA6b02afewbvS1Jsp/HlaVvNpeUZD8kynTS27I
xKYLk3d5V5U5pXGmnxuSzLuxUKp46algX3q+//+awnrp+B9S+JueHS1sDF40LdiqNC+LnKIHHjUJ
GwN8oOEMCdGulpu5nupiM+fER5s5JAykEMDuKkCxeGcxtPYoN4rnU3sjHNy+4yjaU7ja9ZnOMhMG
u4khNr9naQlep8QPRkB0fcA5PwWn3gOruoHthTuQ8g/wy5sZhzTYoc0Ev/uTiy7LuNnUI6vdhvhI
IsLIYpQSukyC7y3wy3sjmWUUcsF/KjvzxTOYQkygqJYtqtwySAk66DcbmQ6E7Ynfp8vpQ6bFULsK
mym9XKihB1EHyQLeUH5gTBppyLIuP86pyLLNe5Y9Ff8jF/viX0Su0cUVdI/eN5BNDGtRaQ/qxi6E
a+Bbd0LIvHokYRPRywRddwvPyCTE+5lfVXZlMV/rOEaPMcekYs9MwE3/jv74KGwPZ9gpd6ywxCQv
eZGAy0mNy2+KB25UdjdtjiegdHKGKEwhqt0cLNvV/CLE2sNS7os9N3DxKbOI9wB/XPzWdI9hYx2E
+r2XXxt7vGZHLenA+QearYxSq33IM9SRdF8sy+A0tsjn9sJEaPbOK5QcS3xwdyn9Jt1va3bPAD0a
KuCbpNhnK9+n3zB88Dwc1u1IU2SB4cS0YEK8fXjHrxusb8wxmnWED8bGWbsBCq5xFwWtKutgx59m
lUhoQBZbAlXLs4ZogfBFxz2YoUfpVwiNyNFOwtvoQcoml4yHtJ+tInERNbYCqv5xSkKzPg/+V621
Kew8/4+iT/spemHm8P+OLDxlk5qLAxIV/TABzWENmGJ4pmXpiYiMJfTn6nvVL1x4AS6fks65RU6Q
QrLpSsMgt3BKEGur8LLoR/OPHOO82/bf8svnzW3AXuytAQR59lJ95blvh1UvkNxCgJu2S9Zf1Nc2
X6coJc9gXKXv2IkiQZmILWzyRpsFgYZNpUwuJpWC0uwZJpblnjSVJ/md0uOTluufJcPV1q3JBAK2
UdHZKY7aNj5704fqs7HeiaSF9g38x+Vc5HmU4dVRvNiwsvlXfRKcim48F52yFz3WlYnPsJknNUZf
W82l3xZ/ltyeKnuwCC2xey0gRQxjXmRlDqfW1sik0xFuNKT5YWikpuuuXtOABt/g2yCnvrFKDt+y
BomJtGLjD5kYtcotISkijbAuG1shAlyzQ+k93pdSTZCFgidA8BmzxQYj/llOSTWNdYxphiXsuOU3
/P4o3vBg9PSGT6DrJtko9xrxkukhl4et2zQhPHXxbs+xziR39gvB8fpiA8EXrjrU2hO5+G0pWvbn
7zD9aj+jCE5YBlmqGDWvx1+IWEDDuehM5EYvb4iFCTi7kEK361VBvn41ejuVjeYNiBruuLlu7DH8
wtySLdcISG4lgjw3LhlSQCRA2O3+c0fWScUwkzvYBPkBtWXw/GqqzH52EqTHG9IXgTjYK+ZQz9qB
YUvAC7gjF660mNWIVoYPsl/ZztVpXIgh9q1z24zzzvPTkViAdNUyuJ31L7hFuB4+73V09bGBzo3u
rsxCyCzSoZUSpo9duuYL1GWkDIoEJ34Kg/kvUPhG5NZDZOAK7fvspoe9XK3+9Ra2Z2knvyJXa6Io
gTE6Pg/23t0IQLCSNypq7hgiMuk4fxsTJg4sUQfnnXLLq3UQYzD6hQSACJlvYsSbey9isx1MmAbH
BvHqY5KYNj0XP8L97iMfenW8l6wz/64wFh+Hn3XdklJRZWVr/rA1P6lWQkciL/Yy5cRxAasCmHlv
6swPF+C0IzaIgO1+ggBkMca/B9FyvGaAsGoUkzpy/nIGmfQVAFrnkb8ErtmZA1sdImTjL6Qm6nW9
vVyLx41QNGfdcYtiV5cC+26/iOAejCnVUQzyI51mZjD1HAswGYf4Xql6apGBszn+8OhWE5VAVUr9
uEA2vCMs6dTYdrPSr1EXkDhowJBM29k3stDITKRZr4ci+t49GkoAPVfn/1bpQApxcHbTekRAuELR
oQtdiJBGXJar/CzLAZ77XIxGZBG91Z9zCNwl91f4pcdL7P3nA8l4J7l5frKvfJX6t9YzbweASMNO
cTwOIb/WNnrhatKK+ckuzXyrbZeMlv+2FWsGX6krmU1HygqDS73GkLKdq5ZcAoOYxjA1EdIQzVs1
6DDidEKsjLuQoWd0HZV6MgyghvSTbJhtCSsnpgqtLy/y0eDIYc4Q4v6XQDiv/SdVpDS5EyiLUblL
DuwWVPsaL/JyszFgQngovvgBZwQDAZCuP+7Pv5Q6Gnhy0ryRERYoqB3RXFBcBhwiDuW9L0iiWnc0
QQcKIkH3LNAqSq2PyF+weAkQVzYsw3Mbxc1feRDALAJFt27SclO2I3bHR7CT1j6rkCAU9X2V7aCj
vyUmPbaHK15GF0X6OmOuiEEuldHVUGVi+o4dquhehpQtcFodtrdqvcNYUbKt6DpMFOescqoV4Beo
wa6Fqac43oeDvdOijkNU7+UrZh06x1cFIPuHq+BNvn+x0oehwKxRJ3H7KimNVCUEXVBIHs6ODjlf
yz3Gq3vjkosBjQ9oUwWqluWnzrVy+G78wLlofhbGMVT0Nv8mSJK5Md/Oe8oz12fD0BejtM05opeh
GOgXWEIaa5MjbAEnAe69z6tvWU0ZFOC6AqZHK2ntTUu/tbLMSHropFPvOyVyw1SZInYmorrbQmcX
w+DNhM2srAyswLFhCiexHmxmRgPF0QQ/TJVpuBNxH/c2YlGFWkbks17PhVtKAHRuxbhLbiu94Oqj
+7xMStJsyLNFDnPQtfUoYMzd83PmExEFVsARy6mSZyrECg57E3d4vDItaP42z4LxI+1/lym6Q8Rv
YLMLKEpove+qIs0hlsbOYa6pxJV3n0OYDmx0oJwx8PctbEKbD6oQvMkwZKdjB3W1Yp3TZWUhmXmo
0dUkJZEpVFlZokri9bprdkN8L1Lrx1ALksAOhcTykEsmksL4Nli9WA3PiSh9OMp9pQXZfgYtcopD
xO8DYoTlvxFJoF/MVlMTKvXiwQWwOSw0WqTAJqMVDHcC6sb3f0mWu792SpOGymC/IcK2pWHntt0p
efUugzDFQeD4uoaAxrFVXFRy46gClKOV00Qoq33L76/uE/uV67mwaziwc2b1WrQyHXr6K1ho23dp
Bhw5gV7HVfKT/yCjM5gBJnCnbNW9HLM1r3ald4HiPoACwEHYWTaIzhxHkxuFTJObGlmm6CeNZZmp
fhQ5Zwyq/MzErMZx3X5rGgAaaa/OBGufPDdqkqusmSgkebXyhEHK7bWKghh2I3NGQjlQhjmxGqwA
WgXTQZuMXJ4k9pCfWYDIXwTMA8n4/Zf/h1/IcYpMH3sDoQlC7UmGMWwpmP+A0P42FwDESF7UgFxN
dll22VdAoS2p3zcAMNR8uQe5OcmCCfhcRmunLp/lKkBeMD+oYsM0t0I7PzUfFH72zt2Yau7kyaa/
MGuvn9kys80ewki60M7NmiHxo7KaHgcZjOX2kH6fOGvnCWhh29DZEG75kLaEQz9BjCYD040VdjNT
NPhFdVngOn0N/gncdZDVUBCnYQjuwQxi4qcEtYuj4Mzmmj3GLxcsHLjc/VcKo9gDRq9XC5vXUkbV
mOQnVinsmHELioMHQkWj1kRSbhIXg6jXf3JUGCiWk4hQIhs8Yc/4EwraWl0k7zySQvBemPpNivDF
sJFoqEnmhWyx8G5cr3r4FUiIBXl0mtJie9+SZKxtNVzUg8dHdchJr7FkrbMpP83StqXdnKNDPiHt
fhs6JZ1qSATy/OzUEnEkDW6XIFFk+wbquNBhZ/WZpybljn0FuSL5x5Gjb7mRppmbEdUX4UdzLn0S
OlUdvZBTac+OiQq8dOOEijciys1gpoVqOO0rs2IQeCSzzUX1VznQK5k/NhkRIXlRM8U8n5N2qMEi
N23gLhOPY8FzHZXnoX1V10+3oRSrKdePPX/f1cH4kM80VNbzEmtTwOmIJ0EzyUvcmZjhMNkkmKHo
M5kEgCbnjPlH+/ig+IFiObkpXc6TU4os6poYpN97rvgAXcdrJmQKAP1IpGSvdO6OQDLbsrv5Tp2o
/VbtTxAAfSmpOayzaUNS4K7NkshaVH5PxqBeS+xh90a7ppQj9ZidpHBLfkfM+oqjs0Lcw4ctDcd7
n+ZzimQEO2OoK2Cgp+zn0ezvnWme1PTIechKhaA47lcI5gTmR7otvfSSixLUoAgMUXUXwlYII9u+
C16raLBr+HIGeNWsCR6FKhHDcFr5N1ULR5lBb+qvgv0onprpHWZ3OJaxmW6nLltqLVLC9Bj4e+fy
Gk1zZ8h7OX665DJe/FBdWVGBxz05P1u7mxXuFTJxyjykhicJ5Nclk5TIXpmuoRes0B6H9yPcMY3D
DfMEBsQP0AMHFKk47uptKNrTWH68oFqQADa8I5ejqmYnjqAtlj8dWKM2XR0ufgTmYBTaXNUeXYHY
bfjfoYQ0WXQox+7n1V/EZVUk0mGrxhRFS96xHt3l0aqmQjAFHtUCZRQfjmSoeRDnKfZQOgHS4m0D
UA+MnXOjhSihRqeASM0gd36ekNFJ6snXQMN32ZOP9YPNGz4sk4vBTXheVfllqs0JaT9lvHhXzco8
kLt4peS9i4A3WfiinJg0LC/QUFakoILn/brgC5Onk+Ljdzf7hQ6QDt1b9mwf5kNJ+1IJVqNjJAcF
il/k/ydOZ0Wb7JZcha4/TtCmAYSocMk2NdDuBrKpuFSHTY4kBbx5+vstdsXgse359Hb7FoM5pzAP
0h+5k7/IuJccb6To5lbACYsI01bg6eGOqepN1fhrzZol6MHQpC9Jt5RtcbddWmjlDLXyFTk3u0EG
o873USMSFuwSxbIzsu5N7brxbOCbcMLpbze7xbwC4hJ7kbW4HSCI0Eax0MWgd7ouWXKgeo9TFc7Y
2vN7eIfm3+faMVOGs4TYEr2RMfbO/mb0ZWy3+A/PFpP7Jz8oSNjG1XW4yySYQ43mA0hooH75Fdhm
l2NblG0nN78RXimPzJe1TZMe0Xw8LUr5leONsr43K0LY37UD3EC3JXmuBbo01jj/QHjQ4gjLIwfr
C6vNsCfDy0Im3bNMyXGDIaDYQWHcoUqadgesDJf9WfzzT0sUa2ScNSUtt3UKtlySprWwmx5Icus7
K0QZJ3hw6Dy+TVLN9jQa60yC+O7vSgwDvkRopBOyBb447CGyhr95/ZKHNAvjsulBemtQ282nNHXN
VSrZLt+3i+WHgXr29pQN/yiWjp2zNn/skhZbRErW5VUbmchAdfVZ3LYPTONeccNAhs2wKSBQmt+x
qdo6m1Vr9e+L5YvbGCJijrvFFXL5bR44MuOPANR6Z3O0SLMF8omzSNtMd3mxEyqqhscHr9oGxHAK
AFpKjRg2364c4gkA/h049tEkAd3ViWRJL8e4tGrCYxW2519e1oQLKSOd3iiJq2hQq6zL8zdffdIS
VLbVDmI1e1+cySJ9o8gZhA71JVJdQ643UmOC3a1Cx5fVYb7WzATSLino4ZuaagEVFbhpEpOSxcI4
0U6D7g8GDWC5R+ArQfAw34QSW4C7+pgVa0qSubOAIVbTQTQmhUsKsf/XvPGoyltNU5ltMjKy4OM3
kWs8FMBtvCWPCrlS5XWeS3p0Qa/igpKg+UxVeDsEbF8Q9xUX/oGxNbNX7sGeVDbbx1oUWChkUwWy
iVUWoEppLMDRMQ7mHItGm7pve2h5+wPoUSEKI4qhTr24Ao4eB+x/+gGbz/BHQytbipFkaERpjnkS
pCFzOUJrp0qHpZ9lC9XjQFdWk0z+P7RvOY3ZX/9kVUAJfFSYxcGUgwjRggBUuGG50p87n0M1bErd
1yw+yQE5kAPeoysSQNO9W3jSVSFJ9YGdqC1m98LFrTfMV5J8vLoU4CwqGYJ66E4ayyMH5SQ/Rz7c
dteP3/c5PoFtY19fnmGetKa829h1arxWUmGmEERxfrG00Hc2OLmuh8DIRwroFXakYQBhfPHtJQDZ
VWrKyycDBPqvC2N3b5xN7+xq+yagJoqV+cLDA0Te3IiiJbkoPswBOh+rZdwM2VO39p0pvGrleiTA
gqpiSe7zYQdDZeH7tK5dNOuXTTxiKbiunLKprMNU4JAmjxS/pB8YXK/ZduY7L1zebXtDD33zOJCj
Xi/d7xoX+oOrFqhZC+z4h6hx0nvEKaIDBJxgRwqPn0Q8Z0lsR0RKLEVdWcMjmLMmdo+ofN0a54Nt
I/3GbLxf4D/rtMUUMW0uBFHQoeZkiioksPzmGzRUeJdhsQlhbWsMfyeCEecMoQQ66fMK/FXnEldh
0zIFj2HgVWK0hiReIkP8QbCo9pvDVkQxK3ESG3Iidh48C4k2+c4q2MwZgsblfiasWDtVFkAajrEl
lUT6Ael4S1PZ6fK3WO2BgzatAkXj7PnCHcNCqXp4m3dBkUN3J8vDNLP5JOTixNKzCHVkbXkG1xX0
RO4463Nt2i/cNMHXGAqd//b63ryrqvsRAEDKojzPb4CofF2kIV0SrTtWZ9fEx7sj3ESfs2ugxEqv
kRcguxLaAQiC9sFIrhupskKPblrp81YEQddCkXI+m7O0wYgbddpxX8RyiID2ZRj7W4/p1h4rf5jk
aj4S4PfBqB8oMhF1ZHtrDAE/ShJMAE8UN80zhjiDM4zLksGX5YV7WPVSomhH65HIVLc8WQUCg58Q
h0/jRaGJTl1+wp0omLV1xU/8yN5w4znKz8LlG5fb7SkUMWZbOAW4sDpd87dwWaI98MuEnlUZ2zhi
OdUcLz5dtqFiggdohYZD6+PJi8NUV6SHREMLwmDsx7sREWVGEL54lSiqYvRCIOhHlHPVZBxdMHkb
bY/VSU+H6aORVEabKOv6mJWMP+qJG4duB3LP1VLIyL8z4VrUy1rWd0ZI6EoXR6WIsBa6Kzr3A+xr
HtIOPxpvDgF+aQWR6DBrZbRQQbGkIPWpOIcH5ou7dy4ZU3G7LNFF1k8ldIETm+eDE2hHNi/cF5dC
yn8mT/eKPDUw0iRVs2Lvjfr7gDYLi0tCuzUQ14dnLpOA5TN1+IzpY0k3nuq/F7uO/e0LWIGemjaQ
Mlwcx4nS20TNsLgXsOPI8rQfmyvIkdWdl62Npqu+Edv4ToyxkBK4QdIJ0q/S2eRD5J80Kx0P9qek
NuPU2rBWqhL53FSI0ns/cq+7jHDXW/+pwKlF6MJVjCYqCMuT0DAuNSoR4unsA2hytu5E46Cd9DHk
ris/FNrEADRcfx5ARbl41+7gkkTj2ezlcbi3xhKdtjzehlNMsojSET0P1XLNA48vmsUI7iTTt2GV
L3hNW7oJMWwyLPHqYmLduhOHPihwwjG9NEWkaSj2zdwOOs/KAlFqJkZ80h2NGIqpsQrVHjKG6t3n
jpkch8wqZTYk7kp+uJL2r4k0U/nlsEJtYoGBAK8IQbN1aBwsu/uU4Mivk9SYzwb5XEcjT4KPPmjV
MgzPEp+IObpuZpdNEKg5TtSN7wx7FRlpWAJu7GnifM9fYmIRRBwRW2WNsKmDl0ywiBibYjefL3pI
InQWcC/bZMJiwV8nT0MWDbkR7fGxcej/DAHaa8VF+jSTTnOWBaJ9z51wPQsYdWmfMndaHKI/T2Mk
fk5VqQMZYtQjUmbtURHXp9WibantLzVvNxtnbI01orSN5UqvdKaw79z6iXes1a3uO09yq5YySZty
L3ENeutcGW7JEKdeWbBmPb0XyBqi5LpSvLqqyhR499KDpy2tASBT/o2DpFfkdwG7QXDfx06Tspy1
W3r3IaBhBJS4QYZfirTDB4jva/EB3UckK2w1T7ompQF1iVk5syzye+5NK9jOHq2E1FVSNxzq+JK+
bTFx7kIL3G83PxK+LWoSWkXiAiElX2FelwLi+gdGo4ANkLkU/PItyYt7GdVPwkSoqr4/yZMf7LJJ
N6X+A1aR45oM0ko8nvGb31mKzOztXI6bZEoge0AdEjGbIClbCEdgrYg6whTZ0QNxW3ib/lgeyjZH
Ikc4RP2oPXxVwc945m7zuFg+ic27Cj6mTY3YCMK2UrFIn8diBmksazdBCdsrjA2zcD8Qhwl1azE+
jNxZBAbHvwG5DFfVFnJaG96IqrdLvzD/o43KNLAjMTG4AfUy7xYWbVzSHWy3ZsfzD51PAKPb0Ohh
bX9u0u72CuRHHz8rMzEITYxu3/9TJUHfNTG4bX9fu2YB+0Qu6j5gACXpNTLfNJpTqi5gSDClUU6n
7K0Avu3GecBjsA98RRNZ/TT9kHSE7k5PpgYTl7b4EOjTupfpOIjeRhzRHJ7hAsK2R9zvkwGVWVQT
JixaGNWGOk9xZALDCNmrIt2EhJc7Hl5R/JuFxXpE2RBW16bWhHZzdeaHU6+mUJtoxF8uDxXza8cX
iuG/CTSYC5mVrDWnW93iyuXk9RKwmGjwcr9vjyxiUujqQxIPJlsAUZvl460YdtVSb+CzeSOjljBL
4BuvKYpgnv04cboQm4icP+zmXQeOVU8Tm69y5L99S68eBRgr5qtr53vfFQK0ZfTynlJN9vn0cpLT
5vgznDoHbgJuIC5lC1MRykmFA0QZ/yYlgcUoNqvv42AaqKgTCs0AUIyEeP88dbPLSjJDmQ2AOHSw
Y+WFZJJdvpnXQ7+VzdqFurPiLM/OTHHdYrW5yOrVEJ/VJHwZEQMfZ4029K2hKfkH8EGhzr7FWXol
D33zbNuJZQ2ndLviEtBODVZSbUTM2bQOJOofjOLUY1jkdp871zWmC714kYN5Nzal1QZPTjupN4lF
N1wQvpO0CZVQkqSF44nmOM3yac5uLvEzp90Gu60sqzJQ2UWHAiysA0nK1SKVwNJkOn+AeNnVPx+P
lY1G6nYBFoXcYiZAoeAJqsMvfdc9Z6egFSduu4bDGC0ZcZTCgLCPqbZvpWLjccCE2bzYcRNs17RV
6yY2jv5R7cesNEKS2y8QyEZoxEjNxbSSjyOGrilJ0hEeUW9zUTX2Q6QzjDjfYp4ArH8tSzsOpEbL
12bwokombqjweCYsX9ZhL8Xo4HoP7pCyMBxpR3BzooFYolDckQOboZgg/ejzootg0DXzRY+p9jNo
WrCis4/pw9XtZ6bHyuRpgvXn83s3KeLFQpQRmuYwsOlBl623HH4M5swEOZmxyE2BVXuJngpXUVkJ
ULgcG23zjqJusuX2FGsruPi0Mf7LXQvkGCKLz84ZF9klXkNE013znTS2Ni5Z/h7+PZd4TK/7njsd
i/pZ/3gY1YeCQTQKzOaHYEEZUsQ/3dtwt8z8yIyG+VuQU8a4kQMSRQNdeNKDiXilmIDeVdFxk7iz
VddyjVvQdhIW5eCuzeIqwasK9zYB/xHXPO5uxcHpevbJq09DH2+005IAbnWQF2kJmT+QbIHGGfCG
xcQXd8s3DZLPARiWzBx0EWbcxkVcrxfbvM3y8daGprtPHWuT5y21dcbkEZGiGCsVrYNfuRb2z104
49tXUJhyOF9dn+xM2+WXG/pPlKraqw42VqjYyXkqRzNLUK6TQRFI5Cw8NnyXrtS/Eud3lKaHnH9p
kwu/qAuBi2s9B0z/jurRnRvFRrkp1o8AcBa+7EjiJM0jJEktJ25KJ+j6eihLUTJIWqKxWoiEgzgz
azxQktCMG+9CynR2UfzxH53VpcJyIHs/l8DNnySo2ChNrBz9VbnD2UT85+tXPFd2uvExx9Lz149X
3wYmsjXKgwKfqtVnRfw+KXQQ1zj7KJ7wzDn7id+TssZ9VJL0hJus4PduQqE2h2ETT5+lhM21JwNY
hKhIGFxJWHaHW05YqtaI9zsySloLsvZsDJSaGlUjNWKB/f6hyd0AmV5eH0R3cXEICjeAwJlB8BT4
e56JVfJHqvFQLMNTewytuoHpbELyzRzgi74cii2Ni8Q7z5hN6MkWT6W+EwSguVCFhbrRsDXse/sn
icD6naVEnAcE+E1uwtmVM7GFhult0pH8TwmtgaRqYkurw7GEFBeJLVYl2dUhxvQWd/dwANXZPPu0
omgG2cs6recaVBLBNDvSKZrWXZ9U85SJADo06h2MTN7W6NaEkyqXRz/3FmaxO/iIJoWdTuWf9V+R
3VMCtoyOTfxwGrIqRIjkzIO74w1BG5+CKh08PUw7WfMz8RCIIm4TyaxqVzAf+BW5XYq0BKH2UhMa
4CwJBtyWtWv8285KZY6XFfodDWDRsq1fgWtGwC2plYNKh6xzmDzv2DNsbgw7eHG13I08IEOHt1lW
Gcbg+cvA0e0dL6rAGLBn9zE5FUXaIiZVt//7hdGAyPwxJbt5JXgRV4T+9yHpizE5J4xefZv5Rora
mWcyV3WSCiyVtqmzZlT4lOunsHO+130bZcAvXZomyEY20HiIp/4K90ML9cB/PlXNvmojSIZFHWDL
RM6X7Yfe2QWuvTf9uHcqxLvCiI9+PIgkrQV6b86DhGX8J7XQmizYMLPS16AWrEBbbDhR6VdiAfqq
vkuev7XlVKzFpavU4UWD/7phD/222Ha5Vhji17I0arSlKJKoynP4z5hjLmPwNbcGPNxzCXSh/bzf
ai5UQbirgixU22+XbPwaYKkYb5h5rpsnDtEg+YfTb2+dBg2/ZR/v/MOCA/fufIvJIOU/rviPYpxh
CZjeKU8zDlBHaZcPRqY4axVOx+I9P28XdTPT2nLCGvJ1SCCabdIel2X5vbY1vcrJLcTFQV4rFTNf
zFdexjo6z6ZU41j1S4uS40TwsKRQcISy6hlfMw3Xn4aeu+wAvEcVlLMot0s0ThiUPfxUpLD0euwQ
cc3/AdOqJHtZdxbOvXPslVpWKifym+F+2ut5A0MDsbrqPezAWscTt82Un96F7P7N8btkogIknCsc
Ahmdos3OVqmP34gVG3SQk80n3CDIdlDbbeIDcjKtfob1frkvttohLk+J7ol0gzgIf4HFJuRVBOvv
m6l3A9dlNWwgsJDeTCUR+AEFpeU0om+dgqLk8Nj/YQzt2Y9J0zCzp4DZLASIHIfrtF8H7O5Q3RcK
J3nloDoUCDvPispp45I3I4zyaQADLHkd5kiwTC1GeCFY1O2140QCTHJ+MIttODsWxKE5TA6/KA7L
sAx5RfbBM3gaQSEpbXA3aVXyjwL8fJTpWGUUnCPSNbz/JAuHAqhMv72wMsQHlRQbKKxREcp2w6Rs
kSIxzL+snQcO6rGiY9GRM5IyIaG9Ylh8IYhIUv0qjFcO5bPyA4l7VuRIdvKUFuCFVprKG1igtUpS
5LYhtkgfKiJtNCQG4SY+1tgnGoMuElBP3eGBwCc2RpCMHzRBlEpTZJns1SBQLyS2uZi1VWUYJJ4Z
BTO2oABNn5ctGWOxBCmtOjpcII9fYHrlYhXJL5HF77GQljFgv3sOX375w3YMNhEJi9LPqNamQjbO
p0hzgqAc5mqy22aCzhipRn7TxWj3OzN/Fu82gGfAP1i0ME+DtOMFwt9sYN0obZiEVGQz8veFBcOo
SuuSdahruYryn/erLawfVUQ4zrEoXN5D3iE/ayk+sKpvIQnFiNhepJLtVFap1oFenDg7ydx2F5vj
vaBRbq8rIJlqz8rjKyGwlZGGJhW+J8HvH8jouhHB9bJB30NgdosQuf6N5UaBqlCGLHst3/sS6pB7
rdoTaJoDOvFGwxNWH3P0i5U2KsmmttdIZW+kG4bha/hKCEDAbFO5S8a0Unfiszuw0HMrEa808EaP
22WK3iC68oSGKZjpr3bGdiNfDe5dvwzffc5YgZGN4wJPjraBL/543fvimas2ZSW0baZuBoohc9zR
VV9F3IKpqaKekoIQgF4nfEGJbsSP6gu4qwlGjX3FotuELJh1LI7n+MO9z50EfklFPpNtuFeyXgtv
jRAnfsSWC1ZY8Z2CrRMjlvr83s2V6yVZ/S5xgqkhfcdTnIpZjCL0YKRCUhG26iJnS/kTDq0rCLcy
9SCYUJkCGWEBFToXCDRwGdL4KZmlqz8ERAlxTKtHXvVjty1knhN4+USfEZXKfPEQjA4kJe+qLg7Z
9WQwUsmn9ernTt+/FMrwfzGciOBWq8DeU9eE6SnTAD8A7fl1YhZTrUnYeFszlDrIhpA4ytnCPh/F
ItuqRNg+P+/pv5R+2zcX9tmh8K7XhYQpV6j/DOX7/npesE/yJiceodjwqjEQryRq+8+5gthDTBZa
5O5HvoV0c1EpaPSBG2Sm8ygH4nl0lqjfaGbp/J2ItXwxZ6S+4i0+Yt9xxF4tZY8bA9IgpL+DBSQK
Vfypnm/K4ZVOFqDyRcdMWN2qAQCvB79MP5gRESGg6W72txZCiaPkexH8/hOEq/uN9tOzHu5Wc/Hx
1E6fARV/Hvw4FrDKatVUc7obilvhg33+NZ7YkO4Bnv/RslyDEwChevZWwxPee7wNt44IJ+ucEwSw
mvq2SBqyZFdh20n9TEjuyARKyZH4eze/uZSY2N/B2pihRf84ccGCGikrJ2Y8B8QeYHyMGDB0i34q
dwfbOmsIJq2ixmSvV1SOoCUTzEQKF813bYbhTif8NY1gcp6BQlpa6i9Lz/Rf54cs+615CbaaalTL
89qYvyd8u0Cn4brw+GNxUzvrZSFOwg3g07RcS3UIixsJljw3a26REZX5RNgHwTFOndCFnUHtvBpV
H2PXDt1U/v7YLG3uGf30rfgPKTmVumHy24L//qnrFkQ6HtedcHW2V8d1EDZLCG7TONGv22r9bgWV
A5HnUU0TIOnPib1x2ZCWc+qm1ZRb2rPfmZVDtHUj+o8rraM6zaif9yCutLmlFP2rXTHkZJb2cD76
XunIzo55K7KpljbbPwbkKSqRZXNHASLWi2oIbAUSM6YlMr71R+cBGHMnuVv5p2fDfLaA5Dn+BJvQ
FRFb4KLbjYdHW4I//cX1JEUAdV61gWE+/3ZpYlT454P/q2rUYJ9/9KvZWvqBI8qbvfY9ck6SfgEz
HHMLkcu/BdCoNtyzwrIVM7ewy1+fcK2BVTiL0Ar80BgRqaj2DKGgbXHOhlguZe8N5aBEbW+fRxv9
iNIY8GxIBE+8KrJTQwCXxwZGNvGiHEtSq4ASTKJfBslU2Hy665jos2DLR5He/ju3FFRUFjcqfmEN
Pv/UbG+ZLC4JmbIs//3NjT4vEBltIsoiVAwKLjX8sxHevUXVmEuLb53flF1/sgpCCFuSul8EYEZt
XI2WPxSbB+SkW/dKZkenY/Dn2WKBsMrCAKPB0P2GaXvqZH8si/ekDwGwOVlL0uxUDT0GKl9Kcx/Y
+UfW5bVx6vOjsHE1cjmxhXBIWPahR5d81dEZkb9UDJrSSi95+GjweqeCj80pS5mYYrHpJNnWBNz2
qwe1CxPtYNaXO7RQ2okLBJ83oqt9YV7FSxAAXUSYBkI9AoqFKKShQZjtgwG45aheeMOjVhVzH+8u
cBz/4vqLjo5QeMJKo5OhQ2RKLpY3hInzWI5FsONVV1srdX+lbUUfbw2pMEauOyEvc7hIflnYs7eM
JTIF4JPPNQVCAItroUECj1Yk8TmLgU+2u7eV75BNzn+D0QEFx2pBBNXMfc5BtM7inFP9YPIRK26Q
Tf9c7xGgqo4UPfRF9Tx0vT+5JmT7e1SS8+ZtHzmHLD0BOS7KqLDZ/L6e+TzdU+nRiic69qZZW9Mu
BmtadusYItceHNvW5xhmflFEg67q2ZVEHZ/MhIqEU5UWVQrR8871ldnd/w7PWcNWUk5dGpXJnuDu
8ylIDm+rMpGZZ1qHkCBpMlxVphyywU6HFgLGFMLqP2Xlnpv46E6ug+VBnVJmnOTfYlonnSFTVTn0
itb4p5f+Roy2hT6FCSPDd++LU5lTDfDigkuBqs9aarMyc44w3tEmvj5M8CkebX7CSOhG/srW1CdQ
es/w2tFCYlTsHlSCzWMTCOLZUBy066XfBeXcJz1crc2fPmGiEWFzq23qBwhUFj7n99F115Cm/CyB
orhtp/BKR/p1sB5hJNExNIbWm74H41EFYA9qkgTbPssOlxwqcUvvYIW/ZZILRXCHPE6iyNMbZSJR
WQHsVMwkc5pWNuUGlNHo+LoA5Z3y9SUVdJNWMvkDfiqQ45Jliu8eXiuoq7phuEv4HxAvVsp/SHve
a6L2GL77GrYNxL+6FuiaB5mEe4sIvj599W9Fptny2IBDQRwRQtEp3QWfUvwp0xGDbwP0WqeiTCEK
ErgMXopmbzlKUko2GDlMsyIcKkK2uExcxH8ExNZm0XaNVivWMw5sRF/BkEag/cn9EbZq/6Lc364w
l+b1X9JnkwtKQBnNES2aOP3uIjgZc8bynQsHPiv6GTrgJDs+F2vG53iHrCH4UvgN5j1r6HHiSVRL
8aB2VZuxwsERaIebBOvJva3s19fLrpAZCacTfKw1IXYqMRlompgOUS7AI4N3lYlAmQAVnqLM2DuU
wT0fQBLw/TnD8IHsr/XceXCwzy4o8AmvHo+ANWrArxj6PpR8O9WAzU4X/yMwCtCRq7aLaDs6hsav
MpzY3QueU7K25jKEH3FT9Ckp8vTjGTKjDNS9XFxmtgAIMPVgge3WZ3JbePS9QSvHJQAl0BlyuNHR
grTpl/solhIyKe5S2uIpEyXGBiDDUxs3KaOOv/bYo8PTnTvEgWF19Q5wlNtVA3wokTrOJTl027Vd
dLDQ+bFVeYvUU9WOE65+u/I5UuGW1/2HoIhe7GYR7FyeOnTGbisBkWNnPWllJdqhezvyog9nElSw
M+Okg36j9TTw/pXRCleNjzeMMFndmXpZSUoq0haf+JvWA/nmg/253sjC2rldMDFPvpflrVvefZAO
3g+1I3ApsAXwkAbgoVTwufAQyE7w2poDhUCNRYVxNvSs1OjiKwNB6210KHlI1LxX2OQ2cJR/YuWg
RCRbEKdSPNodJpercophvsww2Vew/xlupHjmuPkEw8UH4kosKmlAPWVhTexiYwF0K/c7qSxxoNvU
I9WZNRzxuYZ9QWOGeR/6s8yU6Hdy9/w63omyFyMCXAZeSBHcpkFATbm95aGtAl1ef1F5Nojfhbtx
yVCZlVxAAE6xplfJV5dvohkYKt2xZ634o+rCd2edya3/ejvUfkCR3xZg5scXtO01bZQ6fkeDei+D
mwj5BFsn+7vyRySEntc+8LiTEQQPFW/OJSer0rPc+4Wklz0CkO0xYX8HoAV4OAl6uT36R/C5MGy7
51oGj1DFQb3Ss5vJbY9+H6x4L+3ROU+Lu7mb48lPPtzj5DuTlKJbRo6Tc0jHqKMGYsna2zzdus0j
cMpVgi8BRuXRIBD7YhcOlqy4U2uRWza5ast2R72x7MX7Wejr/EqTZaoLKwzEjzvo9RyfMFQLeK8l
cIs1fXbBZl5lyx9j4bStKCkvF+sUk5/rfpgOffjeauXzOAZklKqp0E6DCSl4kK4Wt0xWELdCZOAR
4GcHq2dqYwowpdpSyerFhqjuq8ZDw/Urb7yCewI3Jn+e5HdVzcFn4zYsVR0Hc6B9WUa5UkN0ENjq
IsoI09u8qBipjquI66XkJFmzXwQY5Hmfu/tY0UcUjhtRpqUc2zf+vVmwhsJfNOalegyfQGwWi8sb
P+Q9J27JWqHuYgCnj7USCPR9C35aFuX9FYwoI4edwBXja/LqNnZj87RmvbtkQoExLolUvW6RlQyh
f3UEJJ36QU3Iq3SZX1/VCmRx724l2qXKahJ8LHahn9XWb/EMkFZQy8J69c0TwOpOWD7At5+N13mY
Qr3kRYasdEFxn07pmMKaQlcOTWHR6ZEJsSQoEgbxut9qDKtV1SgQv+CGrQtQSl4P3QIu0O8lQw5x
/R9NOd7fjtAHdbaMmF85ySfp0CZBz1leS3Sw8j7+F5gS3VHdwogAq7JBHl36o8o9eZvbVmkESbmt
puakzk4pisKxnN1K5O+gXvhcPuGcuFMOitp99Mmzk2LLYTOW+8BK41PSApx5yPbblDiLulsZzIUb
LagnDbh4yRPUPdI7BntPovoLVZLUzd86sZi5ltFQswzFrEnp3kVHI9FRJ3hkWhfeT/ODgy1Ll2Dr
LLnyrpgCA6IAfDNzJsRI/TTU0EosBXMnRaxdFIcV/AxkNF31m+CYfN1jJ7VL9iFdQOjUa9KJv7YG
RV1lxoQn4FnpsziEym0OPVlEoS5/EssQP6Ydd2IBvKpW+hfU++L1Med0gqhPjdg5d/p0j52OgjMg
DNlD0CAUQouiaz5bmVcoPZiYHvNBxclqXhtCaL3U4CcCLYV1tNrgXRDPYnGl6GqTRrTaUM3OcFk1
VbuYrP/mikHcApAT2biORDm0pgjYOit0X8V8IcYzFtkQtx2fcv4gMkJrD6H+fYln5yRtFe5L6jfX
gO36ksBf7VB8zAiVwrMuKi4kdE6www64CkLtb8ITzwByXoz4ByameRwG9L66NHATDBS+nerTQLY2
mdMqbbI/GvfJk264Y8bAlEb4xvQoo2VjqUW+WPjFUb05yVdlfPxm+KxkPLEGbkcfK4FgqKHRQCV0
v+5Oa74RuSmxCrZEjUz9E45JY7QZZcU/5tcZYd8Tb53Et/eIhGPcxRalxMxcynQ6QnPMFzXy5tIs
IdQVkBvaa1w3aI7/QrsUFWnFeB5o8Krq8M70WP38mwGW84Mb5g9f1nroDFsMtwsD6GDGbRTAhp9D
87QfPquIoJ9XYKScOLX22GFwfH/6sCibow4EpeKm5VZLBVNMYbuL0e+VNACAtIzbR03286CQs3ny
LiQWB0RmcOMBV8Ywm5BzOcvu13PhPuHeL5J2Zq1HgydmEo5XOMWZHmixTV4GxMaimEgo0yBuYTRB
e2EZWYUSPlQZGDwfpUNIERq5tx8ZEeIu/V6spU1SF9ODyRQaXS5UldfHbYmACQZaJ3xDYhdySFYS
NZdovVRwxvg6/S945QfiuV32924fDD1OWL+QLYKNfVGcJQRmYsQCfGkhpDE2+XfncO8HCFEYLi4V
BjvDt2avqxAHTABrjhb2obU1g4NJpfT6YRn/Sxa61Fa8Cs6yYmE6xR/bAF28kdJD4ejkC2NxSOPs
1Mtn58EqyeW7nvaVw/p6Ymxq9lMiozd/gyyi+okLSA8GrbOEHwG0xapmo/kzBW+fhJ08douQSVsF
pcWeMsqMqHv/p2FwXVUKYW2o52woyo6HCInz9XuwX1oj3F2NxPmwY1xzD6a8pCv/QXzlBJ4RGR2M
1SUziwqHG1Vi37Kwg7gfsKPpsOsTpB/2LLk9W7I1bjtHfzxxvBSwRx2Q4OtV5qCbN3hqJ84yEI+R
Qe08ysm2jXTuMJaqfmwuil+ku5sCl8FvCDi6ihoGx/d3jN2jAveMKvrHHR2rm3dkpZa4uAas97HF
E/DOtGtEUkjXKJ04ZAT7A99VPHP35aaGGLN5DIZOkx20TNKmh3EPP8BVLqKBkqpvw+9ZYXKMp96I
70bGnI3xrtZUGJMzhHUU1vlg8pzC606KV0llEoNcxyjo2wBUU/l0E7PkvNv3iNGBJrevXyd6Vqzo
UIFXjDhEcA3ddHkchua1CWdMRn6o1WD8keZH3NeHul6NFcI/kcrCW7bgF8Y1p13ApCFfo7+JX28a
s34snySzgYlhchmOmEs2rdnylf6Iic2xaBjLcw75NLCniN8JAZRE0aC3LAQQr5gbqPO5COyspH0a
tQYi856yuzdncwmG0sbaqYDeTw7TNihDfR74YV/FeoNFUQe6JgqSit16d+th1aHWxqYmSgS6WEK/
ktQTLeA4bkt3JHbNIey984sleP9fP+9mdVD9wUiay8/54y4K2AbBBiqezcSeLbTOsumpl62f/31F
lLtXIG6mevfmLqLkFSMFcyGzXFMNYU9NqMk4wXt005mxZ++LIVWr/ss6o7h021gzJOS78cGWM6Cp
aXBVS97eYrwch3Z7x5qcTi0RKmWRTUtcdr6tqLEOsKH3/bCSlLHWZachBaXnO7l35taA1Ki/DXf9
84GQY0/9/ZlIt1I5C+EpdSnu4wkQibCVp39f+bP4XhTsEdjW5oT1vfGWYsLvfOzG6h27RudpXijj
Si5x9dyT3UCjECaLzm2Ujsy2IgC9B5D1W4TZde4FOqlDGMa0KSyGKBPzI/OwNZd4ZYJJ9e4SWTaK
0Ds6Ccdlo0v97ptB5nl8u9/jMswga7ISLIgA1OhhNkFHPDuHKZQ8qwtMbj92hQTa118H/JbaeSYq
3dHQiwAvOdBNP3momGnBxmCoSHFbU933CWhCtyEchSceIVEdGtBCVznuLDZjzVykrtzPlLVpLD50
Yh8Hp9Cb7TElm7CRF7HYpDXiRGz/l+QV4mER62YKtwshmcmKW/lYVjyMGwEFs6+PTjk54rrF8vRn
H2Qi41Ex87cjanG28yOHbecSmrzAuu67m+kiVQ3Fz9C/vy9MdvuRfbq2o/s/dQjZYmfuhcCh/Hrv
t2HF7663zMAQSbpazfbC94l3XK8W+PjQExb5jKQ0zJXwB2KherZp7uxQdM/qGeY2pcvB0tJAnUzX
5JJzepRxIZl/aNjHO2d4XUkNZ+KvO+2eVcm94YrXaaXw9IMykNikbS6KDnPNcH4FrDejClAvV/YS
Qpjtf+iZLyYFllYi29EPNSzpjxiMAIuZuwHWRZynEtPYblQgMfYvyE63vItF2MkrwwNCAWbxzd8q
rGrpVykfwtglDDLlq0oGmV9xRDpXRbmddD6dMp3/R7Jg4P/Xv74H1gg62QWVwUja3GhGfmsx+r2L
73NHaao8ysSnW05Sykaw32uFUhSJHH8mkhrqYVSkho1Gx2hWYHGPoNcvqSWNxzM+vbNmp1MmOdNi
Nk9tlB8zfLPKdUBfw+SRewBoItb+eadfkVsYOXV0aE8oZKhTC3h5DOQlPZFxO39UGahkKWvf6atx
xIIbscqn1c9iYiFfx8a0B0FV/fu/oR6xP7ED+rFqBR1QUnbXjwNRY3siwLiGXRA+nvtYzyWGpFIh
kkut62OOHEsic2YRnCpIuqBjQx+gLJnRtpoq7JD5dpp8/JNfePotVGdkXVDPwLdAId67zPjBsR73
mENbc+4TCqcXrFc9KgKQ3JasiglxX/msLERFE/TEoc0oPMKiQHhJScvgOvGfH+ZLCspG76ebyKxz
vv9aa5rSHe1YvpHVBRsVmnX5sxepN2PDLb7exSJWg6+znuJa0ZxC7ZUgwP3uQKgBHKguQjezjx0f
etiQ5aMfHH6vQACMH9I2wMQZ5lva6QJWliH+GRUKFGGm4mN2Ro68OttlOTnarjzCdAcbsh6bnjge
VD4ohs1kuHCUUAApKEOJofi3iEY7qO693n6oUqxi7n3gNMoABgurDi0EvYq2LELN6JfngJ1lByIc
y28WLL2MUgyG7RHWCeEfFnlPLQb0yer/bm549NLpPClns8Et8rokvPIwhblE+3DPvFkEvsFn4w/o
W01HOsgVyyYRLXsYE8IsUVQfsRiiMNwLTugHbeOyCHwxQRlYnlWQ8Q+et/d2I9awLQGISHQodtvI
4nH0Lg33Og2rSy9QrnYoLs35r7GQoTf/9sjVR6/oJBRU/pd8xYHngXk4IVnqAwUt9MOJkWrXY0sX
bXB+EmmBGjob16vpgD0KXSD6YeE/kBtH6zmssjrrb+2OkwG0teiWPVKVl0XwtkAqmLUGopt3Xyvl
IUfIOokmotP1Xe3sA8aAC9f1wb6xc9Atm8fpa5tJqAvKljtgwIRu1OCKL3L8K1KAkrlFctIl7jDc
yULGl8yRrfO5rTBq7JvdobdKqkTHk8Rqs/ePpum9FyxzZraourKb0Z7N/U68mSFRlrseTj52Z+PT
7KBEc3ZV9ShEhzp43U+IGr8UESZRUhX0tZiFbHJU6Pxj0sjhQX4FsQ58Urax5bzKDaXAR150dXXZ
qjbW9YFwtDE8hkuuKH1ilJa8bJGNXUgqhDxIHRvqYuy5hZRTur4VzNUBJEtSZW1TkNJSJm0A0Q0j
gD5fwbKLJwT5xhrcjhz6muQ1RtoKKxmKlf+4Eb0k9RZMNY4DETH2QjMWW18B7b3cUoRNozq7Onfn
xocTgHxVzxtA+z/moYBw4s700ZSzSRGEntAEtx+h/z7I8vvkUz64x5gyPg5tux3sinN+j12dWiDd
/DZE3KxxkSNilARCUyTHe+nttVsi+v0N7l/UhNZ6zW0ofZJupODDXMMjIelTAu+Ci/PiAKmlrRHV
TKmTDrdno8Ey3s5V/pdO4hO6Tj3405UzVSYDxjE42cqsrVCLJRLph/mhtThONtl1WsaiTItZoGr1
e9ziM1OtlH+TKBwC32irQMrAVbUfdL6ugxx0S4EG5r5G9Hu0taQqVH8rlfKcHTvO7HmAtMaFmeLo
LNlCGBzDgHNxddZ3TaiEmWWpeqiGxNjkdKARPUQtYD1N8QykrJidUiTfRRFie9wyt75aB5b6vV2S
iplsocJcvw44nSVVcuNm6R8nCXcLr9M766ScfnB7cCdbRgGLzS9CIcVK7MifKctZ+q6J2m80IyMu
Nvs3+HW9I84hby4+EiG0+XL5d4qFhGhUFXcABuOpIydn8R7gnndsOagjhpWavS0gHcEFPGFk0Z0B
Uhc8YmJIiS3z21CZWaKiqs+UXYAn/+q5UJR0PMkl8JhdvbBTc/FoyFpgF7l14Jtm+9fgOmtdlSZl
BqZ3ESKCqAoOL8lMwPTp7z5H2JHhrbTkLTyXpI8+HplRo+eXnikQTYmFlxEBmCsaNzjgOlL5T5sw
pBVXQCTW+pTBICd+ogMc/HbMcK56KDl5EmStUy6dOtJbk4HVTylONwzaIGjmuNkLD3g0vEXGIOq1
gITuGxWGMMrlDUD5WWCtD6iPP03iB9Zoj0rtjqa7J54JJI6xk3ONAE3J+zm5gg5DryNbRi3cdEMZ
/bxY/F249wmp0bclKAUjqr5bjf15Uue82PGSvahjugcS7F0PQzX88qogDXkDAlFULdE6IuaB0CpL
+Q+OmKFbslXqyob6qOdoUNhIDNsdoPd+O7XNkAnGc1C/qa/CgpRMnSKBgMln8shy+5R+8FJDtuEG
hYIIZ8PX9U7zgMKfSPjqPJlKYnch5LFDRgQffwQ+R11nbu2NVrXq25P7zMGWzz2mZs80v/UxN252
FAENVPCtfB84Iz7N7Iww9qDMg08gWp+0m9vcwSODZ8SzVLklCn5gi9tsc+ksApx8I0H81/lK6CHM
+iyeOzVRChhqlx8VoYkKvxr1i1oACbERue2SuoW/cprHZhvjgPoANDGyIZVxJsS04UmsVNzsbjl1
sWB9ylzZcOSuriYKIkwEtkS7PhleRAxpbQzwWqOLQcHIHD/ksJUx2SxfuLPCejS6jsLvm5X/Z7zS
SFINdfLcBuvM/wuAV9lCwQmYDU/SL+tGy0kKai9ZHZYZDpKt14+n22BtGcFgRdY2hRnMyTiUQUAk
j1KZFRgRdYdz1faf+J5GTsU5laTVkF+TIAvIg0NVNzipVTnc0N1LLv7ib86euiPcOezbcoGKmiHh
SDWl8T9PZQGcrfN/5W9qj8nZaTlrd+6AIZR8F9Gt6eCJg31wwrIg5V/C9a/pShzcPr9ktmgGLFbm
9iHWXch+Ebl8ESKQkNv4dwcPgQQgaWX++k6FpHCq45sJNo9Uhvc+Lv+Z276tiMtBrYVPI45Ss80b
DRq5qwJEkUSxnr16kehYekcG20MsZ/XBB047JQzX8NiAFNWylYhxmJMQhJZOqgEIJIg7leHBJaqf
y597hEbdjNS3HD6AW5mTuvWAvIdQF7Cwg5dMGcX6OtzeRzelVpZCGKP5seeYWumrGzp9C0bJYBz6
N0cRnuUOwVgwd/8GWt5naTn0WqphvCoGWYp3hiFIj159G3cy2UqT4Pq69L0z0F3NAYnh3HfIdC2s
Osy0p8nURUH10r8SDh5QOBXj9OKZvf8UC2O2Scjh+1isi7OcRO8lW1c2k3y/6/mqkSgWkkvqv3vV
kCSfsKw7SK3dQx9HHvmKN5BZH1o57EEBjFcPKCwx102o7htiT2irrKoHeHatfLZfUVNBcRPq5k1F
Pr8248g5TpLW7BDrBTNdNbM7MqEo9/9nKsVmRbV/xKgd962ayPmJAAMIcXXul3W82vqQKc+6+RBf
gw9ks6Oo9rsT19fi3Aoqq2G/4NJx0z/AZxXgFpcYBAIfC2VFWjApjlhSAkaLhqEnV0qCbuWxddqR
v43MRm52M64uE+Iry0ypQig4LuXZdb6oGJdgQ/wNxqB8KSz2AdD0crIBSb9DWc3f1VzomJxX/gxN
Tl56DrPXu7O4lfK4TlKhX6WnMt85b158WdrcYqCs+tlu2bYh3ZJo7HJCMHwtyPlJiA+dOV6YAPRx
q25WcOjNHRMxIHBA6LoJY6E3liSoJKeuSYr4kKi89ZbjHA/4AOHbwcX4SjZDkou8biBHHTl39juT
9FJOln8KQcg/k4eZ3g+gKeIIl/nGpwyt0BR+dPHfIdcncayOZEuX4QVGTuF///ySEWchEoxbt2JZ
ekLtkKpobYd/KATFI5tpM5Jh/7oZn6ybrvZaruo1cEDHOEs8NvGRTDilgtyhZsln8kNTGt8ye1EL
sTgUw3zoYsDY2hRTueFLMCBN4HBb+0cAgEmmd3uxZ7cLywPNL7PwhIUqb9jMgT90w9uhz7q9OqPH
gVTrbMThFETGselfMn7mbbssG5DxSAYpTPi4DgMKGIncBpOU83OU3F3rUBhRhxIMW4zV6aiBgxeI
elsogvNKca0suhlNF0b0lYz6hXW0EEUbTabZlcXkFpO+1gFNnJO4SOQ6R+RTFbguR9/PChew700F
4e+lcpmEmlCAxBd9Q1w15heF1aaz9fEj/4ofZ7MLsFEmzSyBQgNe+MZiLTvsh/TszhbGAgGerXRb
mRtqQ8LLEWWynbG9hGVGM19mk8tOGypY0pwP/HyvkRs1ysLfxzQSAJnen4tPiMGZnrBAq2ErRpoH
TAu2RrkWpiKiLL9/AJ3Oo3ipIoulb2wsZnLlx2s1NJQi7BnBUCHO7Des4IXnoabjHA/cMZtg23Wn
rkfci+TAPU55BB3rRu2T9A4TZ3SkVhwvR0Ltf8j4hp+Qxp6MJ7X4zkqn3NpMu8s6FOEJ8Y+fpSpn
AESHrkkbd5xyWawJOXM3XDOYy8r5bJx5FXICBVqz0/UnKrkL0jlDzFjnO91lTxAPx6mEtYNhn3hz
4mnPdh/WTIPnfG7x/jMOr5UjLTiWw2WjnX8LoZ6bfpL6ig0Xya6v0sGcW75rVRZxBaAdgL/Vp9ak
qCvzkSBvZziTuu5Vtqex0VaWPEFfUvXRWPkAVmQdhPaDR7u8QcBfyHkWn4tqlt5iGmSqgEBhPG00
KKpnGuswae0ZXWXGHILYzgPOm0ua09S8wLixHE1ZROYEZya1w+ig8CRWNHsKH8ygzbPszWr3V3xm
HDqpq6p4UTS6psrwk5b0mDRKeExJzDdc7+ZYRqEnY2V8MJS4gP+Oe/rStvmzSJua0ACZYfBFQJrS
bOiOl0q2VB0LfBCVL5RQMdDwq5u5tW976q3DsIaRIERoFLke2KUeEoVAa5lmCSeRaDIIFrBGT2GF
QxTQ/FGYy8oH6CmfiUBxDOd6i+QHzDjgJf2BSD1yyn7sy2TOqHagyzgByjuFYpSBikssfDsi/+Qh
sVRPxECgyI8DOp5/7jVNSjdNay+rrS4KzbRYfNVSfjZMFAdQ0OzbtDDMsi6BD8toftXPDmsPVhAp
y9V3TOsDoPqnglwia9ZSlkbasb0235tjM0WMXj8hjqDdxJP8gLsEH36T14vfOJ0xQ/zrrb1LVvap
f0u8BMwpd+lRUODgQExAbOSY3Yn+SGrxS+b1nAnkNbZ2ovjGAtrFcNO+5A3wadSVu/27XjbpAHsm
cx+6xnyAhx+083ftIX7XsJJKsq86JaMJmoIM+BUcSO+obhLfZ+KqkKcTMbrWujh5P+Fqklzzms6o
eyEgzQxw5+ShuhL9/1Rpd1UrLmyxj4phZcRCl4Rwy4YIm1SGSI0Vrk6IYvvpyHck4GH+GAeuCpYG
ryL/XQNr8aHhn0+A+f223aKzJDaYoKPklkp5B6MXhcs3ntZGf3fCeQI88fOO4jiJJ0ToWIqG0gSs
Ut9lx86HpjuA35XWGZQK/bLZBlMbnWOEmjtqeGkQXLFKjosI3hRE0NtRx//UgsD6XUtN6P8fn/69
EkaLz8s9XpplZ0xKlJoD561/J3IeZ9bLnToB3qWrFMzHSjqXNu6YqdDX1i+tOSqpSk28+mldbtSf
n77qZFp9MOWrKu8ubkiMyTc4oldyVRDpLBfRZ98+fRnRsQbMjffb3QjtonsueQQv2xp9QUYoTa/4
KFilBQGMTqF+jC7um2Gc5m8oHRymksKPxoNnPo7qfT6Yk/HZZGANKHn54xcnw1J5z1UT5khOQjPL
9QB/zRAJRFD8Er2xxnLrLtmXmbK0TYe6qgigQJDhOfi7sYGiREcyF1VgYacYWrxdSyu0obuQTJ5B
UAuSPvA/1V0BjPJ7EdWJdHqfJm63l701NlZt3r8D1XbrFAOzK9FuCHSnEKGLVO6mfgxZxgq8Ogqq
kqtnJGhcy4LPQM0nnnX7+m19cjbDL1Iy9sMLgNyFiBohbp8Rhpqj4GHoThyiSl62TlYXjevoWoai
/RbODAhLEWsLBYV7J5mmoY9i2uq9DYCFD3noeHeXLWWIbmqMS4+cPpzqwlXRZhNjwavGP3yOCq8x
sSDz+yKhhJgN3fYr9nTe29lp5lITt8CdCYLzxlUgpMQiT0TvKJuGAg5Uxjx75dXruoX6LzvrjhdB
XfIZNTACFsk3qUpaeegg8ofNMJrxYq9iduCqwxJZnDOe6O/kisNaKU/5VxPfGwllBZ7gLsy17LqO
n25YN6sl+vqd0R/rlfN1wGXWpNx9vwv4sVbK+KHKyc2tfyFZmaeGP2ZmCQwGzNUT8ctjGrBX5K1K
0/iBEQ8w+4jBjc5mbAODIzN7xSHkWOF0kvUQL8KnCaVI/45gYruS4GF61YdN0UPi6WFhd8OHDLOh
giNE+z8zMnT+80w6ECuUbbz/bEGQcP3p1HSMkISHRqKeKiHaPLRPz8HheB8Q7CrNxbjhzyhaJdQh
XeXw0PuPdIZJRZ5eFJbdkoARNI9W/62/B+xAlhkBwjwok6EQUPWnmhOOqT3bOTGE2MiHB/HtIf05
w5kk1QHK1+/RJLU+SUMG73xHmbih97HaHtxNQzuSoUGzlGvAlv2pHIjz2WMPMYuj6s3sAsG4yxDE
61dJfAKvBDKJ4MIruyPw2eijni/95DYRcTQROdojoXic+MoiXqGxfO1zVYXRTWGI/pDfbVDbgjPe
9JHsy5Hocx6POV+2gCc5biviQG3Gp+Sew5v8Iqgd7wezlBq0TjUm/E8UbpAZLP1oVzhlvYSmIwSh
ju4X46ZlIh3+m/iqqQGxNcLi+1964ziZl2XNGb3JgAeZmihxThQVx2R5AA/NaOZzH8WVhCqj4nMY
Ivz4YOzqUd2e2MsBbE8S8bnmrqybmLDaGD5BoMuYqSHhKJqOkZ2WGwsSxMI0z6UbfwZxcPyW34r0
gBKevKEdEagu9LzufkPeXpZ2K3jmtwkfCazHnmit/bIf0j5aEpF7rWfrcgtdnj4ogvPwJXhufRWE
XbPgaUd9bfuH1U6jdpB5m0fgjRjoPuFSF2RKxz5zRJ0C1Rqr/LiEDfgOmY2C5jDgwJeVit4wtTJ0
TbRJ1che1xLWiZ7386NEoYWBXO355INpy+VBrL6i+VteSitDgkb1qi1xGumSWTMyGmUCAv8r+reJ
3hXLOkvHBKaDowmjfXwPgCVKzhTXAiZLbHTwv5QV6rJrsq3UwneC72nW0V/4Tr4IuGlXewmyaOJX
WRw5GBoSi88TYZXRvDPCyzv0dVHbo2jH7/hEdK7gqpX6zIw4YcSjs39Xbz58Da37HS4VAmHxHL9z
MhMmdVAoBLZKKGzn+KBssHBiaguaaUUBqJBWH2hvTLohAp9+WpQkvfNvMzTVmAzNCMmrOFANO3LG
XzUYpCl/GhG9w5Ngk9Dbtn3qz+QVy8Lr8DyIR/F9VUkfiay9lzBo2QJ8bNG/cMRl0FaayNd+WUcH
M0V7pJ8To7IJg8yeeOZGN2Xuk2/YMTruEfPAdYGzI/zHJr4fskKqBBAlVZwEFZ8ozRHMUkBl4zHs
qVMZZvTW3YFQp7Zn8t3bzOzUntVqSjWaA1GoZjIwoQHnC8Nqv7g8Xk0AFMHQYSgUugkMe/hPm06h
+0KKy6cJLANwmIUzSh1A3f6DOMXpWDS36OOt9byg4sqMpc1KjHiP2dOVMsVJof0u83q5zLZVpLJP
ijvYBabq4obuSMT2X8iWfwM+JughpcNbs9FZlDCkMvrHTgvlMvmP2tJ+jZ6y2a3QqCgBFI0mUZwJ
UznQnr5ML28ppd9geo3b1BWOok0liCd80+hceicmudcsuzy0DMjRvEB0jegdxplCiSttenQ5s4x6
ocISnD00/lNaHoRVXu9/V67QOnhfxxURUY33eIyYBxWF4LlUpRMdiw7S+gFqbewMHc/EiPEq90Db
H/CzYozXCq89oPh7/vnvOeKKV+uSrjwg7tJOFRwMsCiB0hTUDagLvN8yZIOJJDkXmv316g5BRUGh
pUpPCohtDxXmt3pNTDnIIO/a7Nz//tINioMfEc+3DzLyoN3YwTD3FjpYRIlU8WXDFdpTxmztZn2U
thf3F4n7ra8aQf4bzXoMnSlmZyxcjGHnRx5ZUXMa8QtRa13r613+uJ8Lmn0f9UeGYwCKOLG/vIvM
UcaR/KeRX970bBho6YhJ6puKMIhwdm2b16vhCPUjGrl/jTbk3+KFM5SIrJ/5aWwGMi9mPdFi2V7y
P+w8Qip69wytgE6cTjCRXVY3ljfljxaov8YU+LAxVj0Od39KoAYi1RVCkx4H6618sNul+1cUcsLJ
G4t1jNfF2Fx5aOrpUXY8afOET+uDKTp2PYXEJp88UXz6dlkfIyLenPHlfm96e3WhR+k4Jc5VQTNM
a8WzagQWtqw2CdT7EIbhJYERo6sA0tsVBYlPWOHuqtP7oqal6ennQNQjKKgmCGZW0aMc/CNGFcvb
aPnnWWBI3UhZEdnFAOt6DJFEciryTI/1QKrIVprwlkRTwG0zHSHceOr8wjW7DELQF4wzUf5fY7/1
E/s+8H0GiQ5USU/N78N1bulHatsN5LthUGv2ADiAce9w5GJNzT7T8spv4F0x023CvOQopZAQcRDL
mJgXcD89KTM2OSi3BGgoCCbnG2l+YD5KtIBTq+auGluPwTbAqdnTZiEbGJy5O/xR9WiEG6KUBedH
8yNQNFJiuFA1aE2Vz5m0PlATx+eScsLCy/KEuSaQIStJglVVQUnuzIpHNlMMHqZutWxmOKozoDfX
oeE7xO2K9VKoaqRNLjecyhdEeD67LwHji3XM34QFZt8kWDFt/RZiiCWamuM9blo1i50fM1FHaMAu
wS5/qnlql0uaoAH/CRUW4QUyOjA7uZ76hyy+p5uF4eRTDmgm0pnBfFfoeEZo/UySPGgOcQSpI52W
JwjNi50PyTz6mV/VHBftdfYusifa3+NWmebT9/SFqkhLYbuEJVF1Quuy5i2J4FOtR7NNlwpEHGZ8
Qlc88XKmHQGlKICKMjhg5pRweNFCXkwDz4Afr35J/fBnrfM9xtwbeKG/DuyevSFPvs8sjd9p5Nqk
+Gb28cr1F2pFoaZXN/DDvzkIoTF6SIuKhNGlNU1Wym+6zFr7kkNPRySLosjr3SUUw8bmcFLc8nKp
d04C9Mk0tL8BieDY+Uq0nLl7JnEXXB/uMAeH5+ph1MpkFjdKKwOXK36QW6A5M+lCMLgVhToXNZlH
vi0+byzUSkJUXCZnpkf8IpS14yXhD3UDHAe2SQxaH+aWtOwNhSnmvJWhMwdQdh70sLyXz1Lv7qlw
MnxUbup1Wjk+0uOBHHf8QgktiCeJvz9rLu5cMcisp8yyti/G4V/hM4FPHKrxKLL+KfCtX78kuhHh
xN7BDYkmPHOhPFem5BWd8IIAMb+Khw6XOWxT3rc7hRcc5dwgZrE1NojHMufEr4obsZUEnyCWDthv
PtfPkJxGDKekxj8JnfTF+pUK3+HDU0Pl5fMZd/rccaUp/vX9grmxhSk4DzeLUptc37RccujD35Bz
z7IzcaTMl2diPuMzz79aYLWaT+CzXBbZsuNNDAN/hFpO+m8QdBRnoREzALS7h/AouBAGAZEqQURf
9IN7MmeNsfBohDtiy46DJcE3mTV2t5gIpMIDeUTH/Qx3QS6w6P4QdOTjrxtn5k199FaOf2L0YVdr
hhxm28olC7IfrgHAjiMNXjdm2S86i/x6F5g47DmttI+OsPIAkDAnit1/bKD3esaJAoRyz1ZkrtRP
2lZqHmkK2e09cX7q+m2YtceTM9aKdwXQpzhpKkCFsEQUKPA+dmmvPH4FMUqY1W8fEIPffgADruRN
DhrmhAoTBUOqNv9f5uN5eFzWOAfwLPnJUkJYm3m8OhyB0U/ntDXVRrst7N+4hceg2F+ZU/Vba3bQ
J9J0xq3zfShRaxYO0++C3neinkAdRFlxSmGg2EYDIyWmcclbB/KlRfN37VC7iwfjlrN7mYzUyL93
ELmCKpPnq3pDcy8H77rajDLAAb4bQNcbqWCwoDm8QZB/S8dWHaUoIJs23t8AyB71tzfHTFexkXPX
4fhfWHttsFrBTbJ1SW6WMPjngaHhEz0qc/gszeNVgj/+b+FJdVCwsprUolhGJPDAgpBmG+rD9q0E
fU5CKul7+FDy3TpU80YuRoET6Q94hhYtSx0lM0yhnJ0SJP2Ec2lU9PbvSUI/ZJEbo+T53C5sbwP4
u0InTxE+ylaQE+k8tFzrfQj/J6BFTW74Ud7/DcPWUNneoNDIW2ftJZNbIowUTxHCVR3JMie032OG
VApQM06LO4VbBIHyhKjqZWacjcqdsGaLPWLg7RjZvuvTLib8xcwDfYhu7rHtMU9xRxQLmJ2jiiuX
Px0CuD8xmPrsaEkBIMyFNsAYDoaFpOkI8rEAQF1FnWAXGW3JiU5hhlTSAQksTW06rw1By6gSUhGi
Z/aFLqtFE1HJp9n12bWg0nKbUk/8jK6yNWlGYDDe5DL7o4egRd6ZiwgJRPJZC4AXt4vOc6DWo53p
kZmDkk7Rl2gdtbw4uJMHoD26fXBPNmnMvFQv9YwP+eHTApa3F3h4AETE3q+XvtcCl1Bz5/em3dkw
i6mVM5mposRVdkUn5YJJhBeYG+sx5jw2C1tlkIwgz9MzuRZc0dQDWMVYCBoZ4pVp5aWtyZTwPC6L
XgWd6LETXtcQ6/5IOz6aDVKV1XT6pq/8lLEnNVBWIrvk/aqSzwsctK8aWIpM9NzU+RipfYfTq+QZ
n19/2jyfs6dArS5D5WVyG+wrnrLQ5k9lzGAIzGYx/HVvba0B70dNf4mVL+f9wtaoCl+Y7UPLxJY1
A70+wn4aULkyYekOUU+aN2xiA7uPpDnPtQf1NrQQ7EMR1qoUMlq6zyaI8T4wivmgFLL2PUrTOFEW
spu8UP7CeeBkt+IUlX/uxaETpxqomtMgh73b0xsPFwVULeGLzuJ9CcnYsX8y5JIOdnlltp9KqN+5
7pA+qo4wF3Tcrk4wPcY02gTzMljOSx+G1dEehH4tdC+HfxXtrF+GbM6OKedJEv+czPpyC55gWdRV
lkOu+lOXv8m/TWh/AaFHmGbwVOonwcBWZxbUeg+xm2fjaaPKDh1Hb5NNf//vgiWmSJ/mI/DzpMC8
zz4pTcSSU9i7Hb1NK2EgiDekHxYx2Qn6/+vWbj5obGmS/HXIHZzGPHL+ve3J2ZlbArVAUB46pdpM
rOd/ME5vUwxGs2pQ8rXyxdFQXXf4+bdFDEjLFlKhLDa7jK136XhJc3bgXfddH3cGmSUv/tXMY8aK
/maOhdYr4s/FEO7MkgbLteqRiN211RvjDBO7LpE4kAsn1clRkxMahHhallkv9Z42IblRG/LC1Fz3
R9n50mZmfIm519Ind5U5MFiUogeweXczuGOlRmxU8ZHe/KLMh+mkYN+RnZdQA0r1TxCMl1Py49q9
sVaI9hXrDWj0MRvI20pm+QoIRAISXTc60xO2jBaRcNsL9R4Q8ANsiRTSzBmxWtdDt3psH8QBQyHU
EoPLMvsCEQZ6ldFLU3nJY5Ou65a0qTd/IBX6WFUIIiE3vC3b9PHAefobHxhSiYMKVBfsq6aOd1S/
xXwve6cybedsYxkMRYc3VJL0Pnc93SY4h1CbcO9UHuVWzcDH+LAAX3Ya2CqPCYILwqX3W8M79Mcp
K7od5shRHaaQodqebAW45eF6sNUlTKB1xX4qXbGwj0xzUkVD5qC0vFA9x5hAeq70iwI+6vZjrtTF
eHdLHV+fP/6CS9e4xz6lXoAULDajwLDenxA9pcFZYAmEiLEesMyUqjl3XhCtBhlHzjvN7/ff2YMB
AVFHtiOb8GhVIW3XwY9V7aeXFayEitigEdCsVGvOqPqck4e2bPmP+5pF9D4SKZhZF4uOcqZwU9mw
rDXmGnhL6t2Vrd8i8P9+zc7EEf4pWOefLIOg+kjzTrIbycngjj7an4ESUK50vFt/PBvW5LvVYi1y
latsA+H/tGcSBznPnfR7l9gbFQ5HkN5ioEvQypTAqws9IIh/dMP0ooDKKkT8XhIGvOgDNJVGPgQ6
/nhLjyy8205dhhyACjaks6I4rjA9vAdMDZl5Rrk2lzDUFnnUiZwn6ZncRBjfjpNq9SQouKvZlMns
y4vV1NGpjhth3nVF5Dbrf/nuBaw3NjFZIhFWud3WDd5zKKYi+Xde1P8XCs3NOeeN+ru8N9Ls0Qga
6er3WugvmdNgG/YbWbHrNWVdSdxmUzi2L4YpQRuEUdd+XnNImx1IRAjXuIZ13vhZb/TUZfgrqYGX
k1t7CcWXA1N/+mHld+ylXrT+MLIILBj4ppM0f8r6pIjKLbII1St9OYmt5Vpr/Uqw56iNSggayWqF
KxKq6YhT/xnwtWYSG6JW1qYtFRQX2YXSXVJ47aMUxenABPIMhI5PcKAt5lJimhieUU1U+icJaGex
TXJQrtEK4o8hnBrjAm8D/TeUVbXomlo2m0ExpNUu6f2H+4nAyK0XEziqEVDJqadTllKxiUZnTMwR
KWz6SWp7ojWsq2vAL4m2Pqcu43y2mXJ52EQcDPxvtNEqAOo3J95XhQkoaRh36wPhD3bNooYX3xTM
bTb+2yF7wFVhq/r4vQAkS6wpJPlsEH6qyg3dvfwPNjMfzR0exrKXpwV+9hinRpybbQr710+3uxPx
eQVQl7cUw1JDCHSdShFS7E+I3xpB8tuf2puG3VYTBFQZQobBzfLuT3dM+atdfZTksi9W9pHDBZot
kOy8ZV4/82mDtJ19jgFY7W2HuZRh+CVp0na59k4yD0AqlJTUZV7PVlAZZE42gPc312tl5a9VCNS3
Am5ezVsVXOHqN8toVdEdmDDheGp9tuAy+x3Tt+3YfgiANwCMAN1skHRa4mMi2vmrdrDRHHrTxAYc
eZ4HDW/wAd4ZFg3RLP4wAx9kF35L/+9cQZBtYHVQYiwKVGdDqgi3w8DO/DdsGI08uKbMEiu0qnS1
O/ysvgZa6IVCzLegdEGXZn9vwnjIzuqADBvFwTwR6hnPKvLkZApvyLE+ZZcFmVFbdXGDK2fpyLDG
BAIcnQXGzGsZUd1n+3bt4oIXYmTXILrCcWeqL0prXaXu7oI55hK2TO+ibyjgHiQAlReKTKufFwXf
j1kwxmVoBkfymSmIOXJzbuPlp6KamvvNIcyHACXL0/6UBdudpFQLBP1BG34hwVT8+HGYm3R4fnhk
ujsuUBCh+iC0xc4mKtXtWkUfNU9THGipixcRP4IO3AhHbZ+ujxGY6Kd6RzQHiVO1aLb7T7cop5xW
BfSFf5nNXbB+OmQ2Yei+yaepJeMaw8JLFniCrOf5IhIsm8z/BJn2+eQOnmKN5qxZ7SAmPMD00Kty
/sdyjhX3CrYX3YuMwfSL6oQU46qPI3qICMsI4b6VDwFHNRAqlQXu/l+ybyt0ZLvQmtoX3pAm4fa5
PuU7XJcJaeC4zDw4YEy5N49ftCfRSB3nWOWsRj1N3sNvAivzLfLOAHLB2FHZbh2ujD/35Q+Z5704
VSDM6s/WrCC1f/47hnh2FOPQK2smyyZY9K2VVhMXM0shB5xu899z9ZPX9pkoC7eLeGWEM952daUc
wU5Qj4Wa6Zj0R20sKy7SL9JdTHNUxYXJPWQMzc03hmx8DS8NoZcXJ9xdQQbHPo8of09hMwZGWusQ
R7qSSBCOWT7mHJ19v+LFLcEm8vmnury6pt1d2O8UduNnzVZd+Xfe4JKIvnvWF1IlmkHo/Y5xbEh5
+zgCVr7FnTuj5qQ4Gkh71NeJa8O9tWIXOUxcsqS7WTLtzc5ZW0tjNUH9U5q/n/UREW9tkqwxQ8D1
iX8HiTkksLlMP0gREj1P9NjshqMnxf/XstVPf+zm+j8HL3mO1CRp2VA+WugGtqp6vz/r0PRrghvD
gLFbHv5oCBR8wMMp6dDueKXutRVQ+vCskwTK9M6+0lCwKXgtv3mQVUmFdylLqq+4crv9N9smUg7x
oS7WUxID9SUjBDIPyZJLRGz6eE8qYOQsUDp73mZX8E7lLaYj5kWb5sM7tfS1OJiS+sVxoeKbGuDJ
f5TMYm6KtiTy2pYKx4C6C0w/gPl+IXnfiy1duyX4yjZro/yNRK/0shzz6WZerYTH3Knzv2hqSldQ
6tMTWlpfoswPiJch8904EMeQQcIKeG6kFLglFQO1nFZyaidw862xHtzhc8Ud3U/bSLVyL64Uxvtd
LTCl2fFq0AtLE3kuV/157+sM5DQ8d7r7KTugf8DFIa6lDFjF5vf1qPAlzHad5JfgUo/YU8peRr2S
jCbXZGEpvVBfEiuB397S0eveHro2rZLyl9NoehWo2lh/pIRGG5+vpAouNw7KARnZO5x/2TapiF6E
M2Z+LBhP1YTG0j9j6Yp/fLL6e5bynRTUWRaVIyzm6RTYbxMKmAZw5y4wfOvM51lhO33iC4CMxK8V
cbVih2zCvvRjyj/Z1gnbhV1OBn+T8otURCFwT8WrYd87fNaTYMPh8p19v9H8BPaXsYMRBkyOo1wq
VIDLcu4DGTO1HLqMKzLHfuLjv39Ja5/bYfaMy4LQJORMUatRISwHLTHGLjtU/6AZ5/NPaExwmggq
A8722W92FJCS+0w9lJRh782ckK+ip15LOc0EqcdcLH/crhxLe5/ubvs/4j0jOm5k7bnBOfq8ELLz
/Tv6C0ttF2ubhvSKz9iKv4ic5e4otZDCmsE+wywqXtPys8XQvD8rRa5DVpudPfbMmC6dUC0O6JIJ
FCNqbhMoM3YOxMHD37NGF3x1Qlaap7C9sVJhWkalTZLYfXILiKneGpMJgtlcBQnUXi4IZX65Hiwf
NhEq99ydbCsvW3VOJ4qySZcM/U/vsg5H+2TuUdUkXZ+shtTALjYmzzvv1lbPnHaqGsnjArL8LGPT
9yskBQFYR6wcgt+R3QFdJXJrQ3J2Wm9FAvTAJ41hkmPM4660i/iVtFkXiQXY4xaZhYaHJ6pwEgRd
FUUDBQCTW4k1TVxODo91L4Sh0m5pAOG4Rj/P4dSOF+9SjbAA+ntWpJGk5jhmkLvk2qKurlIz3Wk5
DSRa81C0bguPOeALZG5EpW7ARvG2rLuspriRB1HneHtit+aeCCq4v73YjJ5QgRj7QPxfnvZuURor
upgH7vr70AIDMM4ZWl8I3EowRKpYAgx5DF8JEtwq8OE/M6H2Ey9vzvMGKtamp6kgUwiRTebgzeWi
xrnz5ouAX9tsGL7UhuTd0P3RStRrB0awYeuUaSIVjyqEV2mP8ClTIhGq+aNvVdflS2X1ImE74Q2W
NI2vAZPBdnqWZBsvQvewUum9WTt8W2jy9ZAdghoAacTVojMxkPCvlo7Kx6UBAEvPKb7hmB41IpOz
iSKOB3oa8WRaBZ2cuy6je881d1lLWfow6ezvohveWe474cf29naobAb5G8gF6WFcaxYzm6vGRbxV
kmcJJMJ8QatbwCIT9o3JHuR+M5p6mrVDLDYiZxBBUGatnBdWEdLRLu9OnvzbSoG+K2ZH8335UQw7
UkqmTM3lc3Cm6LZks/B8SfeVdwZXNZvHqacdfafUuPMX1wLDvqf/0dFtqLMD1lRFfikc7bMVzJzF
iIlTJb4vB7tpaBpSzVDS4YCSdQLOuck/d7xq97ZeXC1AwwY7fbzOwiPMH3C2RRateNrUFFAZN6I0
cCelZ3YMxEydrtHsNvDGq08bCByWEVAPJLWXWRYVGvDnmv2hudHPOIoDhVuxBx9DXkYQyeTOEr01
htfm98wFqTsx/qCp6uqfzb+GdKhRjg+rnmQQ22/Yi6YFkCbE+72se3JMmP8TJ+xb0icNyZerqgIp
ByEAIQKhAu4hyM+7SDpaUO6Q/R0LeGM7mkTqOdqb3m31Ns9HkEVJdTBVbRbr+3FJE/uIVOa73OxB
Zgh1pfw2McyGO3juQjGhgaHivSmkyDJqvu8ENmMmSB+weAnGIIycsGDTCrvvL1ji1U6Gp1xU6dmh
sPjuYrqkWvhNrr1lEVtCFj2KDwSdaXQ0pwGH9wppIxYdJ3omID6PvmDLxhHdPj8vuUSX94ihMI9t
MV7OooitQF0+I78D3QjOJUWEGEEtte2wijvGrR8ttoj3gko0CEmi7WVjNn00BbPFFtpW0oFkcg/q
FLQqZmJvZ3Mrnbmy6EzPiLd/5GyH4Keg+tHi4YJDvD1oWPusVUB8feSD89786O78VBciRONjnOHt
RMZe5icf0LSHyLHQSls5Lc5ku0a0iTZ3PFUDAgrl3VwPizbDIkEb23UTpcmd6Tzc0FHAa3bne84O
Gwb8e51R/bJ6REYnQQwTxgv7WDmG7pkHvQUCbAAL1ID5SKNGwOt8jKzlD1JqkfREpPcU2XiWtau4
IQGcpRxBL3DURxJUFFVIG/ZW+mMwGs8CyAjuhtH45a+4ONX/NdCU23QSnr/sW4aVZfMxdCAy/0Xq
sYAI0poSZmD3dzR4iWePewiOz+bNyYDGS4Ol/AdnVgSWqBmiPtWjULAEZ4HrwrkiK3BwfGrN5Lbb
xv53n/AosUr9ZWO/OJx57hIk0b+FFFk95+pynjxhCNWJTF9Jx1eEzHk8LHQjNa590irtPz7grVCj
YYB2EiTV/3xERtMDnVSj7FLPJxH68117tS5wXBq0kZ2GWaeT0+1SWSruZxt5BtAmjpKc2M/UiJpz
ajSRqGAk2GGcvA7dc618qTkmS3i74zDCTEoTfFBfdenhRKONcDlh+3yAzwhOb+STMFvdwADVFsHN
0BgYmwlefh9BPtHfYjWA/XJEZbRf6XBMXMrVIovB7D0BKshYgP0n2bmJZEIAhq8twBnNralp9X57
LCYQ8hBqHqT1LU8wuGP//im98WOKZtH0UEHEx9pcgjCpYoJPHInjHrBWEdoNDTuv0Gw/bndBEkQy
omyF590qCQtaGkdmZGmNaHcZLSn/k9mlU4jB7BV70No6tPVEAHZeGNMuu3vDqmo3WrRyt5r9qeQV
qLMzVYAoXCrr/OEWEpT9GAvNoFUCHUdeBIHk/vySszI6fj2P5X9oqfdN/ZJKmEFOnM9wdJMwWTxu
foeP2QSUB9int+GMILlOMpNMRnq69foJbLE+MZ69B0iXDgp2EXCWuskxUzlin7Ez9pWuo2KKkPGk
pqIPbcYKVGBQ9GIfMV9YF/LiZmqMIHLJbFH99zNpOu7Hkgvu+PXEM3RCfPVEPMRAnSxgChsmDFmI
HRUnU8g8NL7K/EDXsyAKSpmUQyQ4/BNvTZa/AkuB+xXnLX+wD790BP8snRAmEIatFvFmaMWAgPoG
ZwKquwK5vRYPQy8lVugRBIz5aqyh/nk4u38179WL7LlZ9HcVUo8Ai8otEwK/WMbd3IcNCx3Dwyrq
oq6dNmx09UNU0fvqzS6Sb/yEa9pXyAqO7ezeaScpQsum8+fYJqQEoe580kItDlbjdUtpxOPrXtor
uRhlRxRPekxxZABopHPZ2zMM0cPHPi9fzad3sOdr4d/MRn3vFMIEEtb3thmAIsDRG910jnF5vV0F
7azFQLU/X67YCRv37+IWm5Z6dG29dEcY+d+z0x/jQvyR5T3GtDEDLp4lDvAeJtshxaDgCMKzBlxq
akPUvrmUBKXsJtiyj8jtVDgF5IqjO60nFVkg8gVE0OccWwHWvqmu36fs6sGhbiEWLBxt5oj37T95
TiELel7+8Wp4wvf8m8yYrpV0c21WT0tlwbly4G5zlbWVUz+RtaI1piZZGNAdBvwM/eMwysEOj1Mz
xfQ+Ddvy8/Jyra3H4vb2pEptmYzEgYcv72nVyV26oNlDA5tFpnXgrqjchFjh9+TgF9WTEbDdyIXg
QFfzQhYAN/LSM/beeJjgAA1n1/MjV2s/Bot1yZZjskItYMfPVUSdvnb4uZHmTUHQFs+69FHzqdH8
9ANbqYtqdnI+xizK462zF9sS/J17cm0Fo4+DAUTpquXAsUXrCx4eFsBb/mvxm/3UtyNz8e3Twd9X
Mdoa4+3VdyO3WCzZkIkJtkjkuAl1Lu3bqCLNbMmLT0NhtbWTYXr1HamX71Q1VNJ3AYEGb9St/lR+
nPwtktzaSunvJFhzcWLdhMC+t4t7TRY3wexc7uH095W36phPrWpGOC/HsZDvdNkTTkjpuc/nQ+iD
TB71TY+PSx0D0sX17Ls4ssNPkeRn/zUHXWwNl2PxonQy9X7jo2gFFbFz3CxKeaXg6xkXLE+c+M3h
Ds6KwSnoLHWuepAAZAaGkcahCqFItXPn0OdFjNRKulPu1FHvptACnSXyQhfLI2Ps6BpY6pc5LD18
Qqc5vomSCavCn9aG9C57m41jJG1sji+wTpPxOpY7Fz7eIWrrgfIXNU6HJq460phgh2rPIAc+Rvud
Nxu2MzedtpHhmN2qjo1bfwfskhZ9fBpQDr5JN1Rh0rb/HTg94YsAOXQu1qB2CI+jgO3fq5nvVYx1
ioU2mLeeU7QBSXQ0QBLzNiCLQoh2nS/jYmUmcFQb5gZOPVRUv5YBwgPyj/aupP4JB9xvGRViVxra
+2NTFJ4Ua92q1XdEZUmKIbWZGxw6TzPVVUJqEUFGAYQ/6sh7hv6Aeih/TfYvmyV920+6h5eGMY5I
rLYCBXVPdpBUCLNW+CpPyRi2MWJuBFsqC+DLzknyCgsrzQYDIVS8B+e6llzHYaEMAP98doBn+7uw
5FDWTIxId0xJEjNwhKTfMcUB5g+YFfHBwWcduqzdFzieVDLYa4SZUWohwh5CI8ZHNRbtDWHQ/T7o
4CLfaLRGjeRU2o/Rmp+mi3f6Xs1ucHEUMeMohQiNfNoiLuFGvwfrrzHADEbEpMs/pdnLI1GkBTIp
ghdhv61+MPFjeLXgaebP000Z2osnxbHS7l8UAMj78FCZm4SbdmIlfUa0/+SpETDUmim70b0tci0f
qBhbuo/JARpQzNKPrMmNTAjcU4AG3bCO93zhhrE7QAAKOKg3GKhgf5SzNVFgl3Pzr80P3VW1rnza
jtGP47VIuwMH5N0XwFCqYEI74Yc8HRBF5CWShDDbQxsjgDegVp1fMMPontCbJBfjOoQ0fHxyz8SN
bYvNXKzZOh/eRPtpuXBi/LHqy+PtLJpFWY77XBgjleE/mXbX6sNJ9vbAREIeTkSdcadxtMjP6H7c
8hQK2JEC2FzV8qqSl1KL1q0l6NsDqr+qGjhxz6TJX+pxZfY2yLynN4BQvY7rzyU/N/QZL7a0gFZP
kX/AXbR9gEJHkuY/wh1KPWUfdNWF9K1fJ94SpxwQ12v43KuiTI8SoAjis5gRFpJUBuYglMRSkwVw
Z7vM1WF19vRm8xsb3Pno2Yr7oVmlhUn8GY371tRgfaDibsTKIAPxBRuLkIelBaPl9IAP51kvpTd5
OgA2riD2QqBpkIz7A9UhOCCmYEcQ6ATBc/N31B5rKCUEsFwoXVwZEkOiXggwRdqrK/twhhMwpT8g
z7a09PjBItSx7MNW4jKZ9FtFePTZWpNUE7Fc6MKoeDvSyc+U/e8Ub2cMnjnzxSV6WCPf9brc2Vdq
FK+/YoQRWwv89VwTs56/oCxD4Kttca6Pwtocq3dY1xdvJtlF29ZqMCgswcVvJJ0AwfZmhtSHCzvZ
R33YF4YHCc5wQbQTPDegxg3+CDrDqEUpUUt539oDoEr+W/JP35eF1kh4FAN65+R1z9EJvQ+9ZFCh
yAX5ipPy7giIXs5kADB5j4kov8rWMJj26KAimGyMjdmKU/WdaJz14C7VQAEh7WwA/23qyGKGxa2m
DPSXJUsjUrUijrueCEW+uk4tZvQdjdoYb4K64KOWyXfUBYyxQGGNGr6Wyf/Y4QqI0xOW6JwENo4Y
Xd7NpfOgCwQALaQkjvJSII/wnoQkDg3ENmIgKgIxKL2gjUYnDLnRvOTuBaJHOD9jaaGmVgrVtq68
pXhJBjITAiii180iv48AqEtbtivVCzfyCsR1PtAen3GFQczCaxZ7YuFPW/rR+cqpdw5QmpE4x4Zn
ESI16MeAqpNlnzZWTK0c2c/zAyz26VzHaO5b/CrDcOPW6qmvKyvZApAdNye4K5SzP/rjrjRjMcka
jDmHw1d102FzSpaYpRBEcpwWqKBo8hxQgO5ljKqYhHzd/SL++wcKM91pRXGfKt+UN1NqyuTKgOhC
IygtMuu3jz2xF/GyVd55E16EhrMPIuS91jw+m0IEyugcBsB4/NNjtQnPKDJKgsD48J/K/KYaZKA7
n6kZaoAPxica7TFKwgdf0VZYB4WukjAfM7g1zECoL95ovqTK0d8SMGJSFu2p3k5jfF1IaABei8QE
Vj4dF84Z/ttcYzR08WQ8F1DucMaXqZAFA3XzfUJUuoimcb80ov9RfUi4DS75qMy0fQR6XnuKWufN
OcuCC97Muk+eFhEnqjHH5wV8k/dTKG0GMYLON8kYf/N3U5qFz/9psRWrcrie+Ss1Y/e0A/Ie1S+g
aquOBCT5SEzdMh59yf3+9/IXuKEfIWWFyYsBG2hAtOzTfdXvr3umlIaVbJuXhE8vIiO3QQeemQdE
fboWDM6cuAyvYkDySSGlsOopjMvWr/b82dGlaEl+U/w/E3VjiI3LkX38ujw74qeH5UxR8QSw9Wp5
YlfL3wHAM1V0xTB5e6VwdUat59VHIPyFuEZ1ZzT65baqF66vWLeEUGERiclgtfRtgF9goecv/Ofc
HGXcomAAv8nJzWnpFffhjg6Be35Rl41fzgHNd6pf5fIjdWaHtk8MDtzyR4lcwZTdFHUiZE5b35DY
chCb9yhdKQ/2SrQKl+bRQZD/H1uFVLPKtJ13YtZLGBgh8ygdZ7uWoy50X/Or/ucVr0E3cKnO9j2b
G9HjI8x3rnyu5ifR6VyWdIKtzg2g+WALHY48MKuniwn11P8pQvv0UscreBDPk1BVZ2ouv7gYFR3E
dCS1yWc5HeH97RM430deLYN+WL5ZUvhXfm+vUmn78jWx+Lbbyl+nO8vgnInFXCjKUVMUdZRf3IZB
fpDjvODT2GTQ2e2xQj1dgI43wy/QmjQFE1jovMdQwFtNH+opLVOTPJDBjMXakDNSwi3SVw2cuYUn
vM3SjdXJuf4ip0BFLpWNr+tJb+dVksGmox/yeTgxQDbjPpPnfS6z3jLD2swhZopZ6vQgc4v6tF4n
UmT/a8/hiG7lBzrGfFadzGxZ6yDKyw0naNFItrwmD0pnNCc3Y16llt0uqnSgs9PrbSK/Y9IB/NW7
Ywk8zN4RCzeQgy15JjxkehRNZR8SLSfXJL0ad+yyzmdaIu6oyjF7l4eGl+n+g3lpEc1NLrMm7Ae9
PwnEvHfKNNFitC5z8xXq0BmDUl5UNNReFQmIV4kBfsydqnYyYj2H+QhyN4Kwvy/e+/xCiRJzDlEr
w1MznLaECXtl7OBpNbQw9UmgpLI2NQv7DR01TSzshv5Tn1c1hKaN3Hiq+kg0wu+xLl6WjOdqxkJW
DMyMuQAAsrb2kwj/fCU0VqIcIGz5xo0PAwMkZZyxzs4zy69RBAKFAQPu0qxcb6T0j5tdxgCaetE/
sTIRUAGEMhZDpEuAVmR8pMLcv1A6JHU7YxG+hb+IrVAsXAA+pnPDyjKHzlLnxlvZ7PuylDwdfn7w
IqG7EdqZlVkCma5F9pcd8F2t6hqpUOcLVYFLelGBSWfwy4PeryOjv9+plb484DIcBFt4rTyf7sp2
odb7nSiqbEPv891cN78m9of9Ax/st//Iw/lRIKERHtN2hK6+90mQ5aF1hN5K1S88Ml8kiewYzY1Q
B+AjG5PSGR+m+V9aQ7irSySM9AjwfwzPAfM3sYQeggjED3eFxdpMcK491cdiitCmhdS6O06x05u4
e1nM6IKDa3o7qKOdXpi8HW773dgTA2BjZt4OEwQD6veH+VzV2xKRNFyp04awgA9xOenPE8F+mBTJ
nlDhIBFTJyqZlnyYJtG6/yBVSKjE+2IaOAu1E8iYQwqn3ALkLAvcPLR1QVGAyOr9D6K3n0FMQ2Yc
gxKLlAfv+i8mLhefft7tLVYP4bFNXSsu7PokYyvU+82oAYdYx4StnFAb/QCdV3zhdp7UffPKyFBg
nN7NK3BWx5Z5hZXqyjXpEHW8W4+EEhnSJnJ4kTfil+lsVMvDXmWv34lKwHLlTmlnkhfnyab8Xefh
1hsktfw+NN5rGy56dGwpIUpQzlwXWQDT8tabzIRpC19ViCPEpmf4/koT06LkAUE/ggK0ebaJesoz
sCcMHFAkLvdVPKA6pde6Ds0ddlmgbxHaSGwMI2AzzJTOz8R/qN3SPnM10N1CDU2g/wumjzvDu3ns
+EQya7OX8/bMlKHJPrTaON4dwDOTyVOojDlINJyd/9JcNxpPabsDuaMw7SiuJ+Fw9/F9kfcOXnNX
1dfQ+RCqUetmcdPvyN7k116ywM16x266o44yCt0ZD8vfTq6XwTY9kBf5cmUE05iCwTaYQNcrs+cT
eRwVAOAo3EoS417hubxaWsvW15+/Vbhe1Bv9Ip/hbxOVJvL6F/7UTMrZ0HBMIEiv2HcR4uwpywwc
JTBxrBhuWx7XNtHSu0yoO9O4pHuhs/8X65Dd8sQwGx0amYTP+Hp72hammcbFW98bu+P0yMKS7R/o
++RFfgf7WYlCAl6rMahGQDuxH//OjSYEWNZOPo8CHd07nYOGyuqxeCR756XAoFd+h7Pr4AlJNn9o
u9+jVmrodO55O5I7zj6nptdv45iBLgZ7QLWiImuplsCBg/pga0I2iSvPDu1Vt/4czOf8MLcx5/9O
8+jLXpcdVFhVrE3Bw3bGc8nMtATqEQ1q7M+JYG9zNfLBc9yFPfzgleAej+dD2EadUv3Pry/PO8QJ
AesaieIRABLpvhsNWzRyX/GArFxEz7dq94cHEsCj9Nh0tDRjHb/82R+ts9e+gOnXuGev6hpqupGC
Iizrt7epbteoXN+Rh+4HMaCkGpfnovahCorCrPM1E26mvceJgZ0S04Bi4oiBfg34k7XxOgF4iejf
vlfxXrWDqKX4DqJ3bXxBP3+4MWeoHY/PUcTUxzUJjinXeQShBXHg7B8gix+9Jp11vPNcAaxqmioY
IhvUaUUr5xsqm4tpSJA1MpK6HXhM+2J8WTlRYj0pqyLT9pu05kxCDxCbn1goNfkN8ZtJkW5toSIZ
xj7swpxoeOvOW8e0gAFaBIBcjvgMtSNKqSRsxHpzyIgCQLxV92jydT03pZC52jIzHPIKp+HQGjpe
0HC39khwt5kh7TFKUYMntupL4LXcTiFvATyW9HH6noTuRzFDRQHqINXdOQBIwjpGnHbhmF2/bHIE
PVNEOitTzP2vMISo5wU0I5se4AAD1M7/23rbzuBoXvUrL2A3evG+9cTPeYx9Ix9akMQ+tionM6v5
X/31K4Py1bIcXZuWWKyljnoCEDtOaainczqbaEfAneWFHezxV6Q84W4QTny+CG7wiDOQqDBEdI8r
nnQajzstmBlSuNb6irKYmto8tctEy+pNHZtPCwOdcxZdnAL9mj4wfxS6A+ZvW6lauawDAh8UeIjK
lY8+LRrBS7takoTVKNZ3yJhktZeUrVemBg01xA0aLGj/Nj8exehu1OSFXUuLl0oVV2s66XXvy8nR
PXGapQ49505GOMtJsLMvR5eAB2vXoQa/FNhDP68pW2PUKYQOglUVByI112wIXjgHGs21W8SlM/ju
4B3lVBz3QVriI8/sNZmoGWKtzioi6dK/gQ0A9DUlZcW1eZqVwyh/zffcodr4ST0hnQ36P1TOpg+o
RIcXZ0egeJ33OSTm8Ou9qFzOoDpVPhfZWsRIM3So3lTfyyZIGzWrtkBdTz6eDCrHRRAteWlne5X/
s1ASW03qPLzMYNlXs7WinJ7PTB8Q4OzmIcWfmxv7BW8tTlZpFKKfdwAQxT2q/KL1FCIZcarpwDyV
8Wk9wMXwjI0D0ZAMGCV9HTUtB2k7YfuN2Vqr4msN3ce8g0F2G7uB6p3RmAktIVspHjwHGJFRCG3r
Ob5me0c52f9RTfDbWFVQ1MKfi7BvqdIEDbwlJd2rf1wHbVOD33Lr6YSCYy5oMZ62gsI0yn+vTiQ+
m6Q+tp92tqt2WVcO9Ae91FjrcN+GzNRYA8Ve3RncQPkQ19R28wpRnMeoq1Hy5H40sACjk/5pIUxo
+jW8AmOZ6ZOAPb7/VyucTcUgp1a+xGmvJ2BkUKeaQVIaQs9YulFPG/dz9B4Nnn5LYBa32YNXdxwO
6ZcAiZcePrP4AyCDQiEZUyZDDdkIfE2fYB0Msr7n4R9imjaI5518DC0QotnJxkNZ2fgcw4OIvYk0
DNtXchZqA704+/eppAeI6TytUHEozMUCiPuGe+JJqPwl9iOXbE6Wr4mQJRLu50wrz+LrZomYtCX0
ud62t0wRVaahquodpnm+/vMyMleomlWVQ0PLJrkWg858PzF17VWHor/+Y6ti2ypA0+pj5lesuc2U
dmiYEFHxN3mI9HFfh49eXYF5geOn5jiDXVWp/Cjl5SKUo8M0zT25tT5hQysdzNiZDqU79hDIsTAO
wINhyITp53hSnkebZzIgoGUB2a/1lJFsmEtU8EjtqUbOwpc1BhyjC78lFnvsmr+Zr5yZTLwvkVOr
U33DVbD4b/AUvvXH4ZWRcJgqU6RDCiq4t/67GY4hXOZL9IMyKh6D8ZJbkY8FaasuweDSoF7UgR9v
iJN7PtqvDXIkR/00uCnpP8993LOLpU6mzbPrfq9qNqY0YJuAO6+DqE+/RYA4dUKvay5+KG9sHYQu
f/9goeEYvSIQCa3MZHJzjVSldnDpk4G/+SDzzgKuobzopmA1YJhlfaZV20SzYzMGnafxr5nOhYpn
HrXoLvnpIjhiRAE4wVZDSfH6OcChtuMGSTFf0a66NqkRW2nrSP9hHanUYDMD/BPmX85PxN63y5cm
Usz2nscK+Q3t+aa5w0+h9dVePAjRmVt25z1ff3McAZDQoXtuczL4XGXw5aXfcipzuo0JIjmQHHku
v0FzHIrt5GGO2oxwNzz324otTPM80Pa+lOnBueem7++d5JRkcoIC/KMkITAkhqREnj9VZI1Xdz+Y
JyHGvQ+2hB0kNREMZuLZtZsEPSirYj3NI+0ozCdkkeXyKzArS8NJXMBQtrD8MwLYtzsmgDAbNrYE
r7YXCaGLC/RrBXnAnk+alOxwx+HMxb4PANU2RpK+vlE05zYZZLXtfAxH3GVVZD1v01kueuNRecYw
sLig+tbUM3ADJV/TK/lFzPifOj39k4X5mzuwhrZY3WCWpOfKp92mBDncSZDb5U3m2yNsUllK4fVF
CNmZpb0lb/q6pyU1V0nxW/AE99oyamUdsjnhO+vlcJg39eatFjSQeCwRsbT1pnZreExVL+c+N/Ql
kIFbo86AyirOKUNVCEJyXXNShnJmIi3A4a8TTLTZ/TsLD47mdYVJqS3vD1sQN3oPLb2uCAzQK/QD
SU4xl1hH1mX+pZypPNnjM4Lg29n9UoUOo0etBNRxTHLRtmGtjDIGR53Sk/JxiYX+XjLl77usw87D
KXriDtc545585TJHGG8yUkU8mqqpV1rGIlfELEl7EGQrWwe+2bd8SxieSvhNuReDJlDjTXqYJyUg
OOq6Oo2C8pY1cf7k8A6le5kdBlicQmA/bH4VTHJ+L/HRs/hWAo48DnDZHYVizNbUuP10UApwaX08
PYSbeMlcyZUm3KfGu24hRaXE38/6HvTBEdHqljaVbPNoXDFM9ybmU8AYVgFj7rIpbeKg60UHQlVJ
HTKhPMVGS1uOBokeN55VSUB5mT6bIeI03WgYZGsMUz8Cs2eT0yknkSP68EdM07W6J8+06pI01Nvf
ozvDQfV48JdDPEyKe3JmxeOgEiCk/43P+Aqe3LjbpGO6Lt1LfTF+TJsB5g+Q7Gm7KqxmFutBdRP1
soIcVjmB107d4xyxeTI28+d9TraF7K0UewC7yNNq4fdnir+JdYCqFKJ5evLMUGfDcAJrR8mzrZpo
04LPXJomhHzV4tEsrhPsWwB4Q8N0+hO54QjV9F2xg7KbLsF3wFCOqa7106RBBe3hEpwrVY8AYBaK
JBbToiV0GwcFTGmiDQwytr8jzxtk85AthxUcNp2fypAKub1w/E3FXhp2ZHT4h64oRPqdRaE1U/6S
FUGP+ot7j7tOV6SrLbYUFo8mmImZydN6iqR+XXGi48EOJYtUpHmJacUw4HvZU7MSpTdwwtkY4vtD
ZJGZ/sBpDTUlrDUmXvdBH3tFVA4mS6B9vPNvBaNPSzWjkoYXzMHo4LbV2SUDbavQfm1mRkQ5C2y4
S8mK04BQSooIGbtMckDExk68qVEtTV71Qo1G02QcXPM1iAhqhyb31yuOX4GgionplBZF+qKUvQGt
V0HM4dhTVVvtp4wL+DaDco5NBYDkPIiEr0eCLjgSdy+VFti0AT9UiD/55GEdzT1X7HUpAKzjmkPe
qMJ7ovEuMEyG3jOKEYmForolYFztB6bBUDlgKWLAPFuG0HvYmObX4tgrnWD3LeCoFeGJuI0aQz8m
N6DTuVfsszgZSzqhNSjG2y9IjtT/61sHst+J3kKT2hPJmFeX10Ba9oRAwEDyjkCWwtr7Oi2n2bdk
li47RXa2wXBYHhv+Apyyo0SXj6gFbo5Tqdf8UAEcRcTjSro7J19rg+yuGJrlnr0pxv6RwmKwTCkE
DlM66IffFDGn9xaL+k3xmZpElITO96SHQKdkqhV0LrbKlNlNjbXIHr9mY9arix+G3IR5TyHiYqHD
eM1Hfh/ziU5kIhSj5FUsZCulEx7df3Qc1Fqc2ZZ+2dLJw0Ld6c4ej2mrjKha2IX59yYIXhtft498
UTq+hCd9rVpAn+oKj2s2G0r/lXabygdbpKxXHT8shqo7L6du8yeB2Q97qARADfhFAR2IVTaN5qoZ
CuIFc2dDJAXxBrBKXjcPEa1StHJ05ZbW8K8D4POv+T/xIGOKFAVzvMGlqpYn/DSRlDurP1FmevVR
tBYXf2P5qa0k6YNv3xJY6Tw1eG2Cs+hy5n5dBwebyNyo3jDOBo/sqOr8riOpaSRcF+1+u2osgcY8
Sh302ptN8TNM9+mKkVoGenrhpAjgvABWFdmKawvcUjnmdDLfaAP46r4gZSEBDFyTtUDMFIO5hjqR
ExvZt+D0G0rGyklpVgjWvySsqdzxWLTlVTXuxuIsDdo84xnytMvoOunlfHpYtfla2AXnIxxtUwfp
1yt8DjDrz27L8VoGj3XxJuZqTVKi9Ekc12lwB1TDkYt+5YcHuUHziekmscwjbTf7KhmXxjHjT7tm
y/LdaKWs61erHg2lUSPqbG9CKz0zSLx1D27XHJR7QRPLw71KkBFtj91pijhLiAs0naE9YMyiWvNI
iyBDewBoJFpoNDa4UvGtJ4Lw1YrwRBxOy8UeOhj0THfizvYVwqX+TkqJLJdKPjTA+BLAS7RBppNi
INCIoxf7GlX54ZNI32OoWfOvW4tymGHR6XeF/GPLaQHlT8NRnuiWy2W+wzP9MaXi18pQzTFejBqe
6oQ2ArBgG3Ue03Wt/BrOaLrYh7E4tRrh4v7p97Hf1MLQoNAR9zgVXb+8f06rOeqUSAa53OowG1AV
r0XZ0fQtzC6Ax3tx0J3++h+8eu3G6D/TSjvqcCDFeOljIHW9PVgO464OOlAb5dobO/G/uZtEE5Nh
4iCbKKAEmmNOZjhcnhu54uj5LA1etFzQJlrxU6hMBlKpNgGiLVEyDPmQR6eH4BmtExalfcQ2fpfR
IXNhO+v2skK1j8acFJjJ3PMGxLfjPDcfgFhdV406E2Pt/EhEacafinL/CzrsQxtA6obt1K/T2mt1
H0Ao/KEkkny3+RpMwvRMQZxred+sQeO2euIdCNFZjrfuZ7+B2sA3ZSkt1cRZ9p5JRMq14RI8t5Fm
uAhH0lfQe5v+VQEB1vD8WuF2KAHfc0eF0XnDNm2czP+b+uUuva5sLa2EsjVK58f6rQ/nrMqEuw0j
/to+ss1jvXC4IKD3aG5kDvfJwIB04bIImDJGV9oWThdM6nIfu0LvXp/3OIeCM6YQwbc1kCpYNUOE
TkhSNEFs/5fmYQjWNoA/5F+Al62f80/lrrMAsOERIGYJEBuClWIOgmqKsmb1Iw5ICHNcICIoqMNQ
+ENLJ3KXbEPOXH7tCzE9hKnxYaU7rWQfnotvyFexnYkM7dwiNK3bzGQQpx/CeYJ32Sd9Y2QequGJ
jZ2l+zN3c3m0YHQAYX+ZmTujakwJrN4Wc4pWiSLeB0P5UgOAGuIIdlR4/2YNtcKEHdyw/kHBx8FY
nVxgfLsaPowT/RZoI7BOuF30fIl0kgerhTnyl105+x5HJHQJQg0PBII2IJOg3XQOKtK7HtyY69Pw
OX6dO/n55bzL2uQtVnJwnQF2z5Zh75V+er3GeEjIbGv5e8Cvt5BogpmKtlYGnhG0bvdgdh26uVFr
7Cr5oNCt51DoOFy4JuspKKV7qeoc7VytSodDxIL8zkSG/mtLrsc5yPB+L/cxeRRDvRj9PNxW9brj
ZYxsfOPLc3l+rTEd4Juwo/JG+zUjMZByu6kWpn2Ykk+vcF3StJakraB0/j9vmFd1ZCcafzMdApSI
86/pxYG1YK5MDi0gUJwRC4ZGjrP9lj7kjVunzIHfWqp03HGnhL3Psu9GpOF2dLzl150sq0Ul0X3W
ID1qjTPnv9KW5SH55CZHHfSrMkcl3rPWODKCMSWsiZGFdcElE4ij13iEFhehZcCBmSZI28/Z0kQ3
qrXdlCtCJG5tJYoaHvDHBd5KgOGCwK21dp00t6i86rweys12WX5dfEIBZRr5EfTrrpA0obmySlRX
SnGkB7MbDk5f7R8EO3sBq/A8v5VJdYlhvFvdJcTqD+WKQDkCz/aL/aWGsuoJXuDMWKZ7WFwwjJYC
BVp0te2jTpX669c9LsSDHXRufCxSaZ6EoyoehNHsR1PQB4Bw7TyIsv2tjK75deT7b9JdJW+56wcV
jUh0QtmM60boWi0DD4uAYvsHXawqxax4pObR3uEgvBGEClB9Jopp9AHMoEwumP/qbKPeTeEN6/WS
cUScIZrdouC39L4Gi2QVPqn5BcOIIC0xYsRcK6LXX7P6PwEaVqh9HmcM/847lv/QAX5vKq51zgMy
QemRt9A6VEUwzd8QvENnYb6zxKATJYkoSOCNYRuyMXLsRZqT+tWXl5QY6ix7xGuJrdIz7QcAcnT1
ZUfamtZtCkYgXobFpNDPg7U8qZCIaubwvcIzUrziqsx8CEwIVYrwYTkRfuv9DmeN/jvCqsdXgTA8
90cEoRd+LXFXCQ4CyHh72Tgxf8CVD/myytjFJwisYTfdZvwFBeq4fbq/0q45uKdhNPjXWof0gzH7
/RYv88gpYMHmZyTU2k/oSmLSsWwjEnUcfRbco/ErSpLBd/d1Pg31YUEfw+l4d9xBfuaZxQJp9VX7
QxhCMsYS/dmXzooeOiay3yUV1LKdHybFlT4F6r7fSMFMqgilGIjXSMpbMTzRP2YUsGK8kb1b8wou
X+TchzDFYyW+d2wsruTnc6tJxeEARZoywcfXiwtjw8cejaUIgkeDq8D/sPcvyhX20lmC/OgAvSDV
IhZnKj4ZY2++JtaQSoAyd4rQ6bOoIOMTfUZhBlSObedy4qrIlPIHtJ6DHYkXPcmy6H6NQZ8Mk7Gg
cOxazyZgo99rmAvopl3waGrWK9O3eNYnqINu52omybeVZFC6OmS4KKLars0EwmaJGD9CDgrRqem5
QJFTzYNoiToFw+XClmvsM/XBpzDRVBVQ1VALN6MlzK+nygpyVYOlLpYDGbP4gWG+XYe4TjQm7L+D
5NYpGZwCjaJg+en0qsuvwmUWFNbmNfNp1JBdxcgHtY3OQyQ/YX641Lses349lmCklf23eoq0f/wF
UUhlZCRG831wVn0aYtsBiV2v+qXbQoIRZsysIxth3opoEVy19Vyoi95+EXB+CymDj2/0ri7YEbR4
nvxb9mRCNSMsYFbRO+Ud+DNmiFpvI8737Nd5buNjtUl69WVzx6jNdHy/3hLC8aadl32gYbA0qZCj
O3pm5vLt2W5kNond+kvU/iGk06XiOERguTbLzw7oK+fp8TFYRmvjyfdOO4Mz7xuVfjVR9/ATCzee
JoMZNa7xwaXxw/5YeTLlO9cS+Cgl09UoPjSb+adjuU9xXkEPvLT+FUGIP2np7/QDB2+NPfT9GsSo
13yfYGGYOtjnCcE1a912W3lB48i0nQs5M8aZ5Rut3+zQE3nmLtNC9nwrmqaFGkTgqr4E3sThK4yz
1ZJnpdklXkun9LOg0lzzKy+BPKWhd0osCrr/qmEtTsrqcjxUJiY4+r71NkTYZoHn4WJXokfKCAyo
Wl00syhIvMSra3XFH31ZBzlrnfXwqdao4mu4jJQEgzDcoUn22xlBBYImXRtIgx/5i8KPYpX2yNpR
BWpPlpkwlyP+dh+CWh0YUYLI7IJb8uy8BGuVTwI3BJB5xrtySYztuaLqUjyB4VqwzMpkK+d7EtQ0
QPCq2yyyryEpJL/JrgH7TUJMS8ifBg251T0hYu1i/rl3TSakNyGDH+IxjtXrzu4fyUAE5GVcz63x
TbC2uzsyxmDNG+HYFaZWX1X5G4Md1zrQHC0OO2fK/Xh3DBFAhskapzh9yeMPKKn2trlPuzMCyrZF
aS43o9r9ytwUoD5zgVP3Hjh7b65Av2J7/xGtmoiou3MUmC9IAViaeUNyBsqp+9EWmMAKjV30bSXP
tuyqDJsehkbgYW69B5hVQVo59RhpMFXC2y8949KSj0wekcmLtGgnlN9xRjVj1HwmOxPP/dkup1yR
W3Ex3Z8jyrQoYmdtrxewa9xHPLUyt15l7Zs+sTcTu+2cmHMoJifpknTFXjPtP2yjM+CHZFLEEbsy
hGQogxPvF7h8Yn5bqq/01EXdIQrr3Xu1Ahkvm9fYIn2LHhsWbXnfxST3lf/JGqpIXizf8HjtyITK
b3HwuiaFUNhM/B5odlioSKJm0r4TK8lvamO0LUHR1f6lHex7zrTOz4c7QSBld5imcbRWP8NNMLy9
Xvpp8HjkQBfx5zrDUfFbEQ4m/g96w+0fcXdsIdUa1OBu/ZIt5RWdz2ZbTe9RR3dhkj4wD9QUU008
O5S3ECNRxAl0nXsuoaP6eiqRDV0vZg5BgK6C1anDex5zzaYh3785y3BErnJ6cXUyBCRVzXJupHih
J88s5iAwrfuc7tYsWEJtSQ34tsamHTJOqgb9T09i0VGm2Lrzr/wISGFIodux0JpCarYMJR0kxT9g
2CRg8G1YLlszE7S0pf2hh8w1tSOIfzs6PbJTeZsr/rDEPJrUA8TNvabj4vzcPbmAoQlrrqqnI8RH
LhXL3P11HxyGEPdty9X/SJb4vz6XTY3w4x3ALr+sgJnAk6usHW87mvY9PYfY8Ne3MVy4UBTdCcoY
TgDatnSbNfyLV/BmMFkCL27g7ETUgDtgRxOXXwdSh4wZoQHM+LPlxR0USkkFki9K2j2AVBwK93mF
O2722Xu1V/fbSwen2/otVXuY/0VNiRYfq9oCpms5FMnQ8Eh9xIF2J87l0WErUMpkjYUNA4MLGkMR
agmdIMaIkbB43k2NE4Sxc0GyG1jZXFeOsmV2beJWYhrDabI/zzKOHnXEIFIwQqD6uKiGGSsCB1J5
ClqDElGS/cItwpwqveBtAIGzDCtZndgF6EF2eD7Joy2LpAzM3rGQZM+NIfHdLOtTYPtw5J7N6/Zk
3UVwGJwl27Wn8yK6vZcBfa8ORm1Lagr+3hwq8xfSrCjjTCr/tJwaupf6PhAiJwmbyV+E953XnWdo
oGFjn5kri2VdaVBhpuosWuUTAk+yyJUJaFgmRAbl4iUeiEdqRhXT1QyPRLnSaorJ3lst8uWyimOT
wa9Njq+6GG6BEpHFByyYTPD4KtRzAhICb9WDCjm9TI715//OPlUbW+uKu054KvgV30QAcEN3dGHm
9Z+K/3SLd5mfi3vx/1cpFrWo2TNzsbV3Fj2M21QQJnKqG884j+YpCp3aDRlsTgFYVXzpfUQeB8IH
zODODa/YXyqp+4PUqge/ITMWzUq9vtTQ/px0/d2PNv40OQKFN02zPtEzHfJbt1Jnny6uQSD51o0O
yIm4/Zxc1DB67GavkOcsZrYUMt8kQ/W+qRZonBZufUdWdx9ykCckh9i2b0aMmOOMF2ohJ28bl0Ry
/TgwQxWbam1wnikrNRT4bP6Vdr38wHmjX6/4Dan0SyHoTBaCVO450yHn0GKq2pFhS6koy69MHeAT
Nq/SVFwuarV7srrEl2lzDs56mdWxG3h5wNfrX830prXpAcsm31OyZzaYrxdnodmR35J1lKRd2zxE
IqjwqQLeEdK4y3aLcBMS2QSaEO44iHdc+IckKA1+k8f7iMsWXleC8w9Wi2Tkmc3UW6bwD3YVOxKM
osiOKdkp92vx39Hulc6DtOsxg5Y2g7o1E3ixNaWcnvB9EG4HUBo7WLv+fVGUg7XBz1qDGCZcF1t7
o5sIA4/mNvX3HQXfydSl5plRj+SZsRB1o+Hh4pzy5bYBMSh2M82yoax7Xsaw/wpaTy/3YO8DwHlb
X3KaiatmXp1sFIWRNOekJElYO5zCQ7FZ5YRJlIFU8Cfb2ACzfJj1jicSF0W3PPR+/MtnPh6neLne
4x/+H5a21hUsrvDiOWpxpMKno9Gk27ujIz6peu6wBhcWMYrTturA/VBZZVs0vbgPKJm7TJzjHQWn
ulfaI6kPl3CM1eP9QvK7kIbGnH4v/eSBa60R5ZI01ZRaj5rvf4/f2Duv5lnRj1Sk7Qhg7TUpmLQM
zczeX7VwoXItjcCaNvYa+tTP8o8oCdXxcAMMcajobiPqBaoDppvuMQhrTD7M025dJsZqdopydl5F
U77X8ms8FI9CVnheIV8br7AqJi2C385ZR/uj9JDchy4lqz1JHQ4IjX/IFF3G6MB2DjOZZcczSOWt
th0jhcNqxbKLmnL2lGcwwRvgZYFKToW0L5omPZZV5btnrhIkam9kOAvFYecoWXWytqIn05pXR0tn
/ZXnpBEnTRiLaaL3/FInjaC99zbbcRsMpEapHEYTPKVUfiaYFpRQTn+z/zTH9ftjR8hPUh08PAPD
Lh/yjCdKxTrt5L0sdfnMKjMb123Xdlu4vOL0EImUQCMlwD//8AqvlS8d91NKYACsSidHf8c1I5KF
alP5BBp90SEm4+4YPkQo3qst7Q9KqDHBcQAx3zYJn76Q0OQyyakP96HTUXDf+zbn+hb7vnZsAjqK
N+l0S4jap7DAx9TD9hRYXMI00zxoC+2Y602fFiOsLTUZI27AqvYg5edhDJlKkd6nfWw0kgrxBi/s
9sSqntI81y7rv4C+E+uBtOHzbYRzkdXH8WCLWdnWp6BP0p/QQ+Odq7VXy6EmtSQRCYu/CVSDEbhL
IkxMrbzWlCewvzRq1Fa2rVdH9VbGeJk1MqU6vO7mGmoAetmndxLDmiagEaWMS4uHAu1PA5E6zHDx
Yp4QYXTiyqjaA4kaMXRhonf2TVRmwNoXyF9d9/cUYG8KXs5KRmh9FxxL0MP3sHApGCpxHFR42A/b
fq4XxZp4DOpIEjIN2Os9Xr7ArpmqyH5XmKNAgcM3HMCim3cM5fjQJP2Gn9kIkycscGLIssdXkhuV
WwatLus21rtZE/jGbaqbOInDCSLxtpAvmq3CrYmRbRmNzAZI56L3aieh7/kIxH3nIB5Q6454GATd
kLAqAra3xwuSmF7jE7/0+G5UTh4K7q7be52yJibp6UElsnZkUG3A5o1h4sYA/NbhvTxAmV7r1Dha
HQ+JZrsBWQiTLCSg8bnqtqa2JiPvtiC/LS6ZtT8JAHrWlImYTC0pwBeN3bXSohgdOXp4rMV2jkrA
d4mzKG9EkOC70Z88lUcVD6nBQeaNaPH4UQCDKcfFwUzoQ11AdbEJSm3hRWOKm0rl1P3PdOY3562w
/okoAcz70qY3XwZ/Y1IGSYGVKjBG0lRLpclVUdtcP9Nho+gVj4/LXskhCdNoplTd8hJvYvVFzDUZ
gSwI1+1KK+0K8rpgJtH4+XccxcPB9LMBnQwzUco/SbUVAGlFIOXmvhpKl7q47WsdM3Xr5vEQo6L/
f44OimUS0C6E3CjZ3R45tuDe1lFJvZCF6JBj2uAVv7ck6zWWPcIweG4TAC2lpwL+5ZSlrSzaFK9F
8gW/cEPKyESYZC6bhw5VpcgYq2d/fZ3wfxUH6SwCopFyFCJzA3kDVtrt2iJ883aFbqH9VPzNS0YD
wWp8Q+fFjQBBnFK6FTE/NZe4eKuaR8rSy5liLJuIUy3FwwDAufSYWaZsPz0t+cIlwVTCoCDKa7k2
ja3+/14T6wRIiU3RSOCRVjqZ60q7rvwcCicJ6F0XFr6sk2rFokKykIWlrWEEjWv4/l78kMKnM7JO
HJOptLZYeT9i7JFN0FIN23VNpOGIDWGXlqtvOj5ERszQtEdSCKEuXvsFrU+txZfQaSThHnkJC0Wb
MomI56yEZVp6VVFSpBmHM7xu2QmA7CuC9VaWZekyM5vrBD47vy/vu+QCAUFeDfLq0rEi7EMFB6cP
4K46b2o9niFH9kTB5LYj9CEpFDt/PIQL7F4t4oQvvGJKHzXK5IrNTZ8FRbe0SXzC3/ka1/ElO9Qn
kNvDzdo3AMw7/qKsnE9v+TdaHngvWpswO87AM9N+n/Wp2YiG+MJRGIWvHhB7nL0khnnCeDY2gcOR
zy+gkZXL/Yr1PVoTksiajL8JAlvsf6yCHu/BfKDdiClIbolWsir6Xs2G+DqRU2IDLsTDKhanQbjo
wkA+K9U7py9x1ngAer1cKUKg9kytDcHZ3zJgpSiDpgAhb0y6NFvUeTrTylJd3Z/WpV7nf0/GsWqA
K5aa1AyWBUjSRFvRMcSrUXVS1u3UYkYbs95pOc+UVpt5IlLcIpZJFPMPRxsLpRX4rjVlKCm8LA8q
Y0bziJfxWU8ijVfSGuDEYM8tYUbQSXIbiaJlHWCvrtVDU2bSO5GDZVld1ki95wMDl97B6Azts7de
mnjnMYlOvURX/9UQ6PAN88QBWo8aVQKN2w2dgzjaDMlQ739XFhzW8wjJthf/D70TkucRqpyt8jAI
G4NEfyfD4/TT7bI/eFBBQ9RluJA7iP2ik15PQuoL8ubzEKoSqcZqvl6eAUI1nECSU1yTE4TonZj0
AZvrxCym/sZ6TctZHPzTPJI7iw46tlbcibZktFq+ud0i3Vav5HB+VkGgI9AHK1qVTYpJBhTcjp5S
wonCaEMEPLAaBgukmcx8ln0uNZBK13nw30+ZffQtrJjAqoiie85OARQyQBYCJL2Eq+iXq3zzFR9O
2lAbsj2X//snx7w6s9N6vLZuXIFho6qQ0lQcqk0+2WUuIUviuwBbUw5Foi5BmuqnXWgYeF8j35gp
XPLKS2Bdixk0XrwncpuIIzY8GkeAm85OYxTC3XSTiIli2+9x0DYSZBMWFaJRw9REr7UxmBs7FneT
0NO6iXEcsAyQQQt0lv2/BnqCSEbAdPs6mIK45tF5meVN/FGLwyyvqSGPcsr+suXMUgHmdKM9fVUL
omVzxxcghhYJqVhtHyt9czLPwRK28IPNiNhc5S4i8y6Nhnb0Jrisiy8NfkdYP4bidttww6IUEj7X
9cRUGCR0JVyT7+CM0Fs+cZDOwUV7HHOjYCokZJCJWgq7kXeGBtQicuPkLFjYdu5saA+XBZu+2iYA
R12zWQzmd6dDLDq0evyPn6uOrFHfEUtWnXmXFi42+oC4aKxRlX6Ung7xsPJN0yDlYMuvZuJiRkza
JA9LVczFmTyo7h96OexvUOxI7H1YM9XF9W2izhOxTYUQgu2JoWDl171o94T9+3OlygXZbaJZxhd3
qjHPQhpDBFpp12yHm3KegIs1shSAhmSl7z1hZBjz3VnJq/Am3ayHw3QBqMBnj+x/z3Ia7dI6ZJVn
A4DAKJLeguKuqcTRmAh/3nlLS8C9w/Q6z7wQxjXtYBCHSNuBFFmLExaqWYfWrzQtpc13c8O9grGc
gYojaiitcwrHQ0NBzEQ0BX8TVUBIqr3CGnsHDt38raf+7CLiwafEjFX0js5ho9O7pDWor/mrBn0i
E/JWmBJhXUxgEgE26s8JDaEXF6p0CMB7jF4bCB1iVJVktsxaU3oSItF5e2QFXnwblsDNgQvpBLlg
8c8putrkKFbj0/ml6S9Yq/MyRUWdXfSNz2x8EdOrjOxC3IraeY4LD3u4qGezjzHvWHvbbAb7FkDI
lFavZyFVBZJ8snFA/o/5ey49BZXKD9eVOyMtBFdlQSUE2HR775WeS//Lg1ybdxBY6/jYR5CuEOFz
zYwI+wJnj8b5raxg3goap1u84HONpCJLhLFhRG8ILt/EYiIPs1b1KtIt5UcpA3ir3fo+FFC6oSS9
tpPmz4JQL60l72/v3lFaaVNx4W/vnEso4nORpLcL4V/ku2BtU9W2z+aLs5h7wGTnwljFXFCol6Z4
BYNeEUwk3L6nag1INXYAiN0FnTW8V7EjtTKPltgESR1iiVsUzPaOsnhKaMSau9xC7aVggIouZEWx
p6RanBVTbVcfQBRoh1UBNl2WzrnzHR81cCewUvtbkutmWaLnI8F9ILrjh8s2HAUy/nCP7L22jLGi
GT4a9ZNEc8A7EID/PhC453tI0HjZ9zEb/S+0GkcnS3yIxYpiw+gKUw+jZdlGo8yWJw2te7LGyrH4
TCpnpqmduZGK++NSQZBE4wN5a6oimyXsymYr+IFkzIsWd33wnGFLZMBpt6H7KKYStFlsR2fndnKv
SsgW6LHy1HeeBg7BUvXIG2IBPEZE0onds5Hi4PLBGD4wOWQmTsYhQ/9FY0ZtM/kvk/ha6k9dyZbD
xwGKeAaqiJqKR6YZKpGJ06HW7WmMQelXPfHwwJAx2F1m34QFhMCrwRnX3oSaRVsEXzgvTbDnk77h
uXa9zY77VsWiz32L4tqCF2QS0t8tT0kwiTU8XEboLfmzlOpD5Dp/DYVl7mZGnu685G8HQ2o02BOw
FEAGd/NOGUmtxq15RNqaelEBTQpf21fZ0EjfR2g1tEpI7s1jTlAUBzfQsDqKZ6r3vtqIA3mlx+pX
5euPBiDvKIMdZxqZLyq77aBY4PvZYHUA5DOyFOU95ayVHMp/rbLg1V5HnxlHVQYRdfkt4hHhEqbQ
wRg3GudtjkSt/1BpiSEMM8l+4mRynG1hQkIcoqOcg63l4ct77n9Wv5Eb8RtJrzGyyyEFVEk2nWiU
4fhMoUT1eCub2Zhxj76XuXT5B13AJHjj80qeogz7rbuW03XLhAKUFpDZtkDWMkiyG5tBlJRZvPZT
bVeyQDxCSJSbdla/lP95pj4+DRVRByDB93UHRF5QPuUrEa8Uje4L8C1LI1LWaqanvWExgwTOucT7
RLFrdj2sEAsZzExQVlggqNF844MyBtRQZ83rWNwS7pwJe/f+SV4d219ZN1IhSXysRQkPE6JbYqiv
SXm6lpYF0QpygvbAzo1eJCzLRrcqJ4jfk8kH5KenMh7bTk878FFIWRsuSslQzoJVrcmEcaOfpFnR
Zgm8Ol+aIaVn0/rAE0gvUci8FNGaxj+N8cZM15PDWs7CaOVuTSC801MonN6bfH5ZjroaWHwRLx5a
sjer5VJ3Y1HrSC9wShUFEUcyFz6rCv/zQdIxXahKtK4A+QCA8rVVFM28GB11nYYXg7x996j91WjY
qJ7MZzo7/Gk1VQQGTUMrS5fL4js39IH6HPkt58C2pNDjhJwMTspx+Ke0sVEXOInaeiR60tYykZuv
fCcEZ475ht3abJD0O+OhEYOGei/28gMojq8uN3LHyFr0nOD2F6gZc/naWhnHo2sC8c+DwUJNxeNu
gZ/q0XbWgFasNlz7/ogK8DqUFBVk/cvcadbhLkcWoabymG85TT6REkNRqVVw/y62KNxtdKDY7yb7
6coSOCo/1AAh1K+T3rxONK87kippTo8uzFznm1fYEXo+AgBhuX930o9KdH2j2LmGOP3wsERScaJF
dZw7jTE/mCufNoCK2Qb7cxLvsgdAcUxD1w28iVHCZbohnviRrGwvJtmZdgUGkgXJlWZBrssBKsSb
H3eVxKPbweQAsUvlMgvCN7IX8isRTbkpL8uJzNzVEd7xyg8VhuYwDD8mOeM0Ga3wnagvM562AxQZ
KNwx9plkzlK0mvYbiMs3JEvUYvaBR87x4CkpKaSP7x+/CYzoq4geLq1mRncttHqvEfjQwo49cevQ
HPCgoLpqh1SjkFVe7ciNLevOCfhceTC4Eg1zPDHSiwkRIVCa3tMXbhpOO5g0ge0gfsORBpbdGiXm
hwy82Dq1WYvQAig4BsY8nAPIerWjgh0sEnjAOfJJL+NDiCHlYs/1VoiYDcGtsPo1IgqnL0IHUBSI
S3qoCa23qNWsH7fDpi/F3FR0foogG4hSpVDYpHYMDvyaIt/pI/7Jp05896WBqEl78LpkO6rQmtOK
KpA4kF4fHt/gbep3MUe6mWFvtPLzFJ09/ZkmIaD9VmKTII+K5lrK9kQOkjnVBIr0F+XeQIWgjf+v
vO/su215Ia7O4SRuu8BTWAgEzZrMVyFsPo7ftl2TReWlZooTK0vfiwH41f2AbgObVlR+q/on1L+L
BYT9t80jmYZBY3DGnjJnuvYap1aGJyhtbeHNC9+JwITRa6o4fmQUZIOrFD1A9RrNmDOkcLAANTAk
qJOf5ZPG40fUMqHHzILOkt0SFwrpmffcNxHUd/jU0T4z2AU6xFQnrpHJbj1c8bwcjB6uu0z2ziGs
riLIzDl9e00/BpNhpWwimyXREcs2eMl52FA8bsCSeKN/MrS5/9HnebfhWn48iHe5luMxWqvX8Xde
5+d0KUgIvrYNMg/zZkWfqJ81uk9DLajYcPL3MTuZyYTrjxhP9qmGinbicBo8XiPRH25W9zO4DJs1
8vKKeS1SvI0rbyugY0mo37TKqNU+55KU7/5DDpEs+EidnWwFWeI+UMJcPJ4KPZ0NFoutdWz365Qx
UL64f7fWE3XXc5kEHiFh6puU0oH8ajgAo/s5New99/qcNuoe5pkdzwcqs2CD9Zsm0g9Dh5n/OpGk
a9MyeGsjX3KQAOQJf0gSzm+uDuUKAqtByWx4l20mZiCm+19Es+QEG5zLrbvu2+eqUcf5CGwbP3JS
waRybH2PJnChjltiwC+IGtrvCluNJ9KGOc1g8yBpfN4nR3efOSwb+lpZB9nUVi2tGGG9vCDuI36Y
UEuQ9/OcUOOP7dd8eGFopWfHEclDYtDhdFBAu8X4VbgUo8qUQMtjKCVpmHwwkASHSPbZGW05xIB7
nY9ZhJdvs7sz35xKlQmobKAofz3v3Ltcy4k3oHUl+Zj8Zxcgq064GHDOlts5FU+c7PWYl9zMOS01
hDRyg55QqxC54PuYJOjgipaDvTAItptDGBoxK/P/sEhzLeP4T7OxxE2vuczEmcgpqBe/d/w2toMK
/kht4YpW525dHJtiJDA40pO4KqrxHCC7YqB1WNCP/00E7SwpZmc2BlVietYcmJ+ljzESHg54RCYv
vcFVA7wwynESkPW0vrB7lznClo8B28GYmr3byolfu4BbuMxi/gryO0ZxJHh+5WSJXNKzVyMsMlh8
GrQJ9IgUIC9s/QyPplzBWvekKotFcAHa19OefMH2swXEzfqts7pON+qQqxnlIWCA4b9E7THENEMI
gjwfMk3MdocifaMKKqjVchG/NTUqKMJeEkX/2zgT8FvrdVdiDLDdVFvXmL6qRKon3a5iAvxdrOmb
7q9yKcyIrRG5z5U1UWWRMdywjOqywzph2ZB4S7LxlvkNCMXom+I8x+s2l7JNX4LvHTFlqy+7faPi
1kNCc6HHAEdlfhTn6rmTGxSDj1ZPPopCk4oXXwbwkAgETQ/eQ4yqB9eiqaVuiAN7mZl2OF72gjYr
KUgIZrGKn/q5cwDXkfTLeNYWNX6g3OXfbTGN4yHy+927y/wGfrB9kyFM56qx7dquZubpEHogYrHG
gBIJvKt7SyrlrVqgDh9G3gOswZMBtbEq5wQJGDxKjXAPSsth8iBFu9YtEhfdpU3mZIqcp7cDSlIf
UiP3DwY+uq6FbHMt/x3dOwxZWhcM4D+9zlF+4tnLroiHfU1r/AdpMUYjJzooQ8eq6POnqWUh/tea
oJoOT9aBtOWKHopsPbmqM96rHWWMxP2EKFeqkxWG3FDs4s6nbytVPAPmtlSkPxmUZNWKL67xIlBs
z2B9eGkpa71Ck95ja9NexUoDBCPRGcM2D55rA1n9esa/OS0fowKo+DZbEiLnclUAVXMp+qG5B0z9
Goju5I8qXFiWDAiPqBLFI6/QLFXo3SZxNKWrf8Rv0yATFRJMCE5QAHGYdJItZq6NQdvJxm3TZi/l
A9aFyG6jthxE4scChIpVjl73I2+wHOW0FWuI/0OiW/dmP9s/9cGJsE05qLxTrYs5r1LVAL93qwZq
6khwXjkXd/JoEwqjjaX+XrvtIKRFEMfibNKFjwGxYuOzPi4DwTfWSZK/IokUx8Uwq82GILBzbrum
VmxkOoXFytuKqMfYwRsoZ2DDQIpW7njmMHK3RPkmL5oivyKMY96D0ARZTgJHjxDRpiE8JBHX0u1N
lhf6vKmwrys1LOdZdmYruTEj12L/Zd2AedgOn94VSgUGi7EocxWI4RCSp0Ljlm24pYrqRlRdXVgx
DT+hKkk89kTLKZNuL+WVK+TwXiQJT1yGd2Xbj/CkmJ6Idi+cINxjBongHZ3BDVsCAG2oc1xgYmH2
acxndCLD0tdJz2QnBfBC3WBkIz1wwW/jxj8D7GWh/lgSzoIvU+Y6InQIiC0KL8MG5rCs4m4/HDFk
ZERFLvK7Z08WJKZkeJPmPZ0M3L3PtaiWDAk83yeYrDUQ484+X2vA7xoUAcpKdh/B1ufxN7iK0Up0
bAXhf6SNcIgyBo0rcx9I5AWjhUPdQsN+/GMmJRIPkoQB7YKuMDL2A+vz5O/OBw8dqOvW/oNb60Wh
UUsz25i8RxZzaAZM41FVWrA/+rKkcfT4uM+ton6HxLstSIi5DtKevs3xXdZtAeT4NZA7BmCBnatq
Ab3NXJcFh30Ta7hQuQybP3rkBP/96YMaJ7QGcehdDNVuyklqw2ZaON3TMFNTpMdZmjUyHTcNCMlO
+dXrIMeVVVbxgR3qU4Hb1EjaBQ/22p0rAI0Cou5CE4W20nTVUZKF3LakU/6hr5Rekdf89/qHzASl
5VD1aNKYR2/8kuwI4aTtvSAhkQed9XNntnP5yph4u/aNgLOL6on1dG6G6pNVEjMtV1BBPmRAcCLk
r/3UZD/T2d2JFSmVQ9WfKkQGf9zOvMmU5SVkaPTrochEFbwhZmCwCbt19UvzocDgX0KuOouund6V
FqtOM4tmZNBvW7gCfpp6hjPVlrD/dXb6DtzUpBjnC4ZiuybzYsRBONPSAWxIc2/BGhe0ltKSyi4+
uTZkNk/2Be8LuoXv2pidFt2O32BHiRd6MhHjtQDRq2BG3MSkSVnv+4GS8Yu025aqVnuP/xSqPGzH
ct3Widkidin8KRPYNT8Bv5OyAXuxuIt1USoEoHUbedxcHJtr9huvyXjAZKfsVaOCYCMWeW6knh+C
YgMs3tBerfAZM5GHJzL+HbvaUBPNcmpxYg2HjxwHIJwb4k224x/HfZu/7v2pcWWOUzVHzh0kLlBY
PuXwmFvxJ+oZdBTLDVhxM+Z+0WFEZ4ilvKlKxFCu9W/qXnOUpI8skadM/WUZy3+I2Y/IEOLv6shr
6w6PA/GMgPxxnrCUVVWBJAO2huVzV6nCQkv7ldfWgiBxVVnlGbsqC+M7KaiQ0/VUxir+wbJl3Z1R
XVo4/QncW31unZltQBFeHwmH3UjwVfLaRJU3lX5pkH2xU6Di+0ZzB7Q+1TlGTzs33+r5Y36niaf/
g/++rGjM4VK/i4oq5JkvRLFg2YkouAeqRggpC/Vgzl0TsGX58DErcFCi+gbwV1L1eVxTHmS7HeZj
dLGXlSZB+JDVsow2zmUDbyIuI01wIguyeee19lZhJVuqdxLNUM0IifpebGYvaxnRN23fpHdKI9PK
JsgJHupAtFPqp9exHrJmB47sD7ONUDHH/7Du/oXxm+girrL0/5MrTOfm4JWeBWda1H3o2MFvHkeo
Jywz8BgVRVBpJ8/bXi2ZqvsW6zMHF1vTNIXrl2hbwV2LqbiI0fFYv8Mu9dKeu5Fw2z6SDswkesHR
dj7g6BspySpWlZQMdSqiOqeyb6/zJawORTeht/PFjdodlAwGWh9/RI0HBfiOaFtwaveSI55IxypJ
tEYOd4msHB1IYRYkJcxLCtRJ8W2ObcP8QlHvS2ypk0o0V8P3V+AOhJ2C84qVqgnkgZ585pL9g4ZL
AAfk/b2i6XTYyc5ERqLsq1+B7zN0aix0HnOcpYas7e4o6YTmgsMSbhaUXWrOoWVDYdl8+NoWC5Pt
D0ZiZIpMeOk9qCGqNtsRSOjhe2bQ3Qwl5na/SHy8b0CoZtIbGn/diWRo0soITqL1cvqmqlQ/57Ep
3pa6qAAltFO+QkGFjiV8iUAeOy5Pr+43BTb4iYqQr3laNWd3qsBa11+1fHNQWU6UUT5+hwzEMBdA
nRPE1Mawk22lV6TeeVeXORXtioS/iPML5lGqR4f5k9ez8iCUDGMQIJtiU+WpCJNplSWGf1RuhYsP
I1gGrOvJcP7ugv5mhS06yS95fbT0iCVYf/rX0DgdxOGNQO/6/6L0WHSUoRNzxj1WOw96QT3bamR+
NsHRzQgzo/z+IkqmbPpptUtpGwPOYAUS7S65I9+0mI2SGEiVAsI9lG/0Nv71QXtZMeJp3zDDJ9B6
VP/PVlTOnxxj3s3XeCg8FWk4XCLh8WmnZGMk8NDv2WAEhcdhmjIBTOsNkpEtNbfS52lXuQFmg58v
r1z1FzhLecrTC5JsikJGHauMcxC78pFxntg4u1UEkXTWK+tRTt6F0Dye7KuKF9Eb6JL61t0CK/78
p8ayZrfYz3LN7zKfdS3+vhunS5dkvwgQG0VxwSfY+FE2KXUACk9BJ4zqXH9KNb/jdFWuWcJD0hh7
SLWzxnA5xIkkqERvhTfeNjMOuxlhmxugKlIIZMySpEG5Zq6c7xKgzi6+i/4tv6pI3FhS0MtXDJAX
ERA71ejzqMbhGJZTD/B5w6sOx0uRkn9N7ellJN7Wd3jYCQHV2cbp4a5OX5SBQpyutTSdUeaVfhIA
phSQgNnLImOt5JSPaPWtPp+/QalkNy19WgmTw4yth0d3TKV6NUavJopvPxxdYAKD3kIuDKe7Yt+J
RuBPw64MIXuUjqKdnkkoNwL0LX1GTKS35vZWbzkJqQE2Fgdxzo58k10bNhxHv1YlwouhKquoCgv9
gY6UN2gp0Apj3iuJLFtnUBzpQj+4pzUSIBt6O0RoCzxoJJxNyXS8lj/Mt2T3Yu8bacoosjN+2Tc5
+LprLwQmMUCMCi/Icpzt4gJ7KH4oUZl7J8kKj0u/MiLhznjuTpnSH2nGf0aB0PZK0MztZ9d2EyaE
XFIiB/DBX1UAx4YD+NZNYtTADhDKnBRSKwrrbp7KjDMoweC4XkAQzN3EH/02ObH+BKMjsrYTgCCY
q2s53NZJ/9y9GRrwwmhrs7FLyT8aHJUfQETq+OkC0JxMSgTbRLJPuK6xzHPQ6F0tZ1K3povKvhX5
9VexiJS3P+FWHbtSlCDwbv1ivZ9bi2IjdCYUMew5PUAuUnk+xsx0HWxRBrFEprh7/lZCwNWahMtb
2c0A3AlR53a0BRKKBaoeJgzjD5OzH8fZ2E25ep/YIV3SS6IGD5J2V9vxZeJ19929hZWFMTbu9G4Z
ebHZvaGDqr1T2+dsiaArZR0KigOiR/7HUBaC1sHlzzc5Py9k+k5MjH/vUgWTLMAezA6Shw5jntjC
jmRedWosR2SfGIfWwcAQw9VqYil+RVUyDKzZ8/KtelQiw0vwONjAmNMCoeLXcjjC/7LMsvgT0WwB
qq8pMTp+WzMWYDiUZpUjg51aEmvlPoIrTTMAJRDDPT/1bX9v9XDHnmLfT/cPrx40rO1o2qFZRpDj
yloRVp1v+E+GX9scnEFPJIqiZeZAUSPEOvKLZ5MphM7qhEvXmcFgHspHT/hrAycoOMUi4xxKFMPM
f0corQXrevyfS9V6z1e8qbTzgpUeo56kdOSXB0KElqaDNMXURX7E/0Rm92+Cote0qvLjuePGi6ZQ
b56vc5Men+FDhz43ub1J3IUfVPOO0twRhlBOJB4nEthMvleYhHWfP8Y7B7M/zOP/SIYeCUqbt7iN
CKiRRtPUVYpxPslaH9KhVhu22ZQS2WmRlrab9YPDaOvEnhfb0vUtrOmqHq8cc63bA8NEOinZy5ew
LASgL0nNlY+xGQDipJvNcUOKUpbOkIu5VD5cGETVfhZIB4SBYNmOzXCSCU1IODwdop3zydJ70r5B
p1d1itxxRBK/b3MmD+WBuHovNzJ6/hK185DL6bLWSX+qKDpCBLXli5D3UmjLflemt7CXrFghm549
mpiTi/2Nm7QCZOvPWyqRGtYDKMroKw4nEZmn5tFVWOqHcwq3bS/B+pp/8J8M7onQ94K9mb+7gYz4
U4Z/MljD1g2aLL/sD4DHcuSdzLlcmLvVO9zzlerO5dIp/TjEmvpbKteuotUm1hGWRR466XIVICie
inPHs6godidpH+g4MdtpoROFB65cZuzL5VdTVPQ1HaVBqAi8V4zibBVNwWH5ZikKySoMj9LKJMXu
UYrBcMFpnejtdoWfG8dNza1KzlmJK8LRNTL2bK/Vr/bBuIqqNMcK0N2mgr171ikF+hWObZUhSDDJ
Mt6a7sagZeDvxPGbOZjNTkr3tpPLXZcQd63U+kAE0HYnYxMwJso94o1wKsRW9Gk66uimklNGIU5Q
ivy4oCf/AAiehcgEMkMNGUHPE2w1sJZecKQX3c7cTmAMLl6tskhl3YNEN+0Z3e97UBcnMbkq5nZX
BT6VFmWH3WK1k/BaP/kE3s1YAcURu3iTuyfEbnAuWnYcK413GzxL+Ol65epSQCLnLitHazMT8r61
bBj/MhkCueELYH5j8CkthHH5jynBlZUfB7LRcdavdEa6GCVsVqgauvgXek1Fl3tkIcfL/siSYvrt
ogkPcCk2l00EwRvDguMnMhkdfHzIOH2iHI8McWlQDs6+DLXxHB4iRX4BWsx9VEgx2jTizl5BRjFh
9C9sVenutPyJlGzzl3as7gj6nYI1rrrD0byXA8t0j0B2TvYj6ykxe2GrhEt/ba4gFSCtw6REDhFS
Y/8BMqm0ce7i6Vd8OPYEV0gWTRd6/P2+tfVODyHJvs8oB5Nk7/pJ+anuZr7ToDYR3QHETtoJiCG8
A3ZUtsAAlC20y0C4a9Jt+An8fNFEGZMhVaIXdunOzwKRcOkrjLTNYa9v1VEwS0HCvldswbww/FxX
kJTO+k9fX7haKer9CLvWWT1q7RWA94mVdo4Cx6ELBPVi2Js094UOVTe6Wls0P0oHstgqn9UdG5RQ
N8HFXTQ1iE6IapPJKalnoGPynkWvFcueMD5A9lswnyJJLgH28IN51nyCdjtsHJeiHVdsMmaJTCq+
DW8jsGa/0qxC8yPi7WWPiS2AVoahwlxzNxolDYKwZsgCexsAmBxwqAjWkpNYyE1CScNnDgS1W8GZ
jesCaJcLN+NFwEdlxKL+t8OKzc+n8fi5Cd7ugbL+PqYyQYSH3MGlVEJerXcKJ+RhIJpawYE7GpD2
oP0NROA6TrHD+gkQOBLTWr5AzolGtehr8TaGfNDWSJS1lGrHgqQ/8a+oD8SkFbVE1eeKNBsDUxLG
GkDYqZ3ivFRnBNP3cGZ+o6DU+Geqht9uDqfSX7gXVLXhnZBiaKj6Mb23J254AzuqK9RpILXvrPa0
F/1UPr+h4xJc7Rm1cVqqY7tVRmiWXgYi0AqPIDQx6wf+JVnP8wuXeu1kdY2GqAUhuNk+IT4MwXJM
vRNemdE6zeHYSP/xwGxcS7M8hIKYGq3q2FEOzVmMc8EgTS0jzmioLKBxPMNqSDxERvXeOV3r9L7d
pNqC+t2XduEHpMbUD9Y/ndv+fBrTrVL8p6Dpm06/6P76e5nO59zncsd68fwc+qzpssr4WEl/X2Qx
5Rzb1qVc5mwHCjFHEvbe05AiVpoCYACakFiBYV5R5e3qwCqlaQe3TvjyW1gfnUYu7RjgAxDhPfMB
daHLNI1MjV0QJQQrSJ3GB19TKH0d1Juw9wT/gPr07zzJA0UPY/aXZfNCt9oC2r/SlytvIKp6ArhR
U2PRfY7iAtyloOef2piuMUwPQ2kWvxpXm74z5n3sTOSwPMS90OHADXxN0gAnVTPaw9HVO0UBaMBE
gxdFZ3P7zSI0m++uXmHCJokzSPvb+hzcNyft2liD2fYdgKsW0BZGnsIbUPT4FlyzOKWNa2D3ZtLj
7tbCnr5SUL4eHo+jLydllRgvEDNRD/3vO2gYpyx8vpCh1IAvMkkF49CJsTJwkMb9VpB0Km/ESYl6
QCin0KngNSU1+2jQjADp4JuJE+WKir341ELnPDxIj5DGeag0cQo+UFBXcREB8urYvXKCJKvp8Wka
a7dfS7SjWGhTj1atc5LrRFgD1+vTbbrEu5czdDiXh68/6agd+/nZs5aKcuXxODReU68UhNa9N9Fo
tkJoTGZkZWu24p0WUvMhm8zkL8QrVZGSaj5VCLhtLbuhBAS1rRP4F+5MmCA9y5kb2ZIgQz65Fd8W
Fs3Y3OnwpZVoZLmOLkq8k7hkEs7+n2gP8RYGsZ8Uv3v1cDNCGweDNjaQN3+1nN4wiWvu6/oZ2dag
zBCG2e7uAFWw/G/8Syl5FdKp3QJCL+83BiW4Z3/8bZTEhht2i4+IuhoL5ZNeU21Z5Pkt1bcz+33+
SysHgSKjN8oSrZpfSJPIJCxBMSZk93353Eqs/1AY5oUBy7FA3KUvGrIrHKPk1IEZMxSZ4xe2lBy6
dUO2tzTXW7s2eIBtEJf0xvX0/4Ibb968fonExmo7t42eQg6TzcGGTopTOlXEQe1wrnvcDTEEwO+9
DU7kSFZTT5uj7t1VbrN8vuR/uHEztmbVS513EStJSvphy8Wd9Kxc+eVMMpLZCEk6V6GxH/SOWGkm
2/ZgufNqqltvyOJAUK3EsJ7nQR4OFmbBXp02IqZ91s+YfsbKQ9YJtkqRZs7sxiE8XZJhb+5d3inW
e96VBCYJGOPggHQ3Vkkc/zhFqnDbRfztcdP6HKBg4QNkfbWz+Xe2z+xa0vk8J4eXOoaPVpSMp5UW
XtzGcb75hEzdQFR98NSWIc7T1NnOwDSRdVJMm2K7sO8x1Hbzbo7cB3MMj10zVQrd3jGIOoKuX8xg
ckhDlZDwv5S83zBaaXeLFUtaG9GHX+0OiDJRmKUTWWpGDi5h/0pihfYVNpFoJRpdPf0wWQ4e1uuV
J4dhIi6ZVZ6/vnog+4yLEEJTm0HPRR3hkEMCDTY/OOpHmC9eu/3lXH9k4XBa/XhlR4DTSAGfCE9v
3y+hDjUIIdNwxe88Arg+ZFZNvD5NteknXK4F4uvilyKHgFBx9qMlbKhFNDcLZUw9c+7hk4vGqcXg
itc5z/P7y2hfpZixlup4aYPFt1PToGD7+fnJzjitXryp++llkx4EPJlfs+s07VCEUuiPKJGJBoiv
UYQ0uRA1AQhqBd2rIFLozrogBboZsRvJWbNAmeF77DDuuQVdVsbqizubX8rcTL3+OQFiHhmIei2i
XGrAHo0SRGC2X/ijFHlSdnDRG6nZMuGPBffIzQnbK5cct8XawaX0bkE/qMM6DIIjE0YOj/Sl4GHp
hHN0EdtdXvPNvp+u8GNhekMBwoPY7FegdyKXRbHVAn/j0ZWyoURBPZVRGNniiTxhiksL3JtID4tp
m4vsHZh9rAx7l5tNaCbdQGgVvGeYBmTcw1DhGeY/g3JV0AEpmVjPVURQsGZ63pDhYp/BykvI5rHa
rDo+dEUuPCP+0nTvwPpggBeW+L46v8bORhJzmMf/5rwZY5Dl5AePW3fDNZU7scknc7UKrx+D4DDR
05R97iTr8WNfQIO99KCvwPjVbA1Mc1twhNf6jRI9K1oL4NXtB7XityLPT+OQ/CB08UDwEkPYcSLt
1RUfIzJCfq6vvS0wYNvj9X0vv4tFgo9R9IbM5YEuPvkVWmOWFwULGouiMTTKTxy6vM9Aj159F5an
loF2jmBXJ64EUnxUEhDES+Zpl7rCLzkoRgVF5PuOuYDlKItIW9FfgKlo6E1P/uwoqv0CMCQwSrmR
WyAk2YF96CUmdFBYuORXX0AFIEjRvUSjAC5V8wY2gKTvW2U2eF9gJo+vf5C+P1FdfH4RRrNgLZ5k
j8MuEhkWIRna2hocb4kW5kmonYZNFmwAMJ3lOwCAx0hrNG6EVOieljfDQ3tCkXn2eWg+Tn8fk8uu
5t1k7bgf7T1bUU8YbvnmaC8Am797G7BUgZ3RWzIY/1SQwL6lL6lCEJRa/XxsAfkbAuVkRPZV+M/A
59bRgixiBdiFDTizEZ/Ud1TMdVD1VIu6bM+1qLo0ed4yVddMJblfBHoE72+IvOjPwRBa3VPi1Crf
4FYJlLw9q2bWvpq0wZsrniOoj3+sCFQgAK6gwdNZN6h8Oj6bOAnuCyfhNzel7dt8Ixhvsa5ck/tD
Q5/s34ll7hQTuRtuVlbYL0kEfSojbAYqZ7C7KbUCwKPCmSCLY/pPUP4tVd5OHbghpBBPkDQlPwlo
g7G/MkOrVfyD3PTcciZeSAMzpgWwFqX7wGeWXLbUNyNZbkRWcC29DWbu0GmjjNXjWuwJP2xu401j
ciK0umD6zjzw63eiNDnJAeIX22rx1xtlJIUSRpoK0yfRZTnTTgN2oY+kXqFapofcDw8eCwWODU6T
Fki3fONuXPOASV1n/00d3Knxg8hEHrFsJCxN6PxifBfblk2A5ZbbasgC/YMiQuZE5ZlCM+puj3A0
D47NzmecB0oF3qjrHoPiq/qVGmB+XEIz1b+NSDxVpwOQmBd9JN/bywfojrICHBA8V+nAN3Fi3iRz
YD+1cQehwK9Dm5skRoRExu1mFM3Cggj3p8DDR692+rz0BJ8ycO1eNcrvJeu3stk7angWUFwCANBh
hVINn9rA2dLJ2vYOJPjiFCa9Dzpv4ItnBloJSTi8bvlvHyC9V0fDDQyNqYGOWqqvQP2bcnQrVayg
IVuIa087q6PDVdmb872J/C+87xMgGnClyuq3SNZyy0rQ65RvK4EhuIbK+AiVmSncYtUaevLSVArX
o8M60FtxhZahOk+XpX2NpTKPRhZQRZhZHvK42urdD1Y3akm6jU5CWfqf7oYyg42Thgshk4tpsghp
5MStbPttAUXfVAh6Eljavx0HyjzJRqNkAVzt8amQay3FeqL/nN3LlBkeikoFT80VIL6PPoMd6mXe
UR8GmNJVHOTn/9MNaKn0SDJK1ctad5ulTsL7Uc2rq4pZaOICPMGSmVjSm6HSthnx3jVAeNyn1uAL
RX6m4yjguKD4e372ahYq5XwlCILLnBxpa4NWxi809xvCxKfwSN1EwhgEkrZyJa/Qo8kti7yYxp1M
+tXLVJWqoM57sXQRsBMTX5GX5bElQGdbCswU7pCaxpFbVVH7ZR9aKZXvGMxWTdpG3w5m0Pvr/zJh
Bm6afv4MpGLENEl1FTssCPE7wYoUMno8dS51qhFe2ZVGctF5T5p2OqFqbQPvcjSxZpbBkHmDZLeQ
Xgd8pWDq8xXyAQYCKtubE7aaVXK8Rzmw3zx2sRJIm5ce6x2/8d4Ew/vnDPV3ypGL2cB9bO8RtraR
CpXdHtOmd2zhIh3bpCmSj6aev1N/vSf1RdZ4EbroYd6ebIFiTCT2Or6ahw/QJnJJBjpvBZuaj1H5
yXuIyD0YvGFDFfw/VXRtq7n+8hakUKlsAhgP9wH/Uno7Qn7l8SSPnuhhGd0rtruTZe3t6lVIpSUE
CBXfjMPmVBUr0o6LMMMhFk5CQHAy4pSApy3DCncKez322ZJlR5EJyq5XdXzh9hp+ccmPoh+PEqzY
f3E02Vy8qmFg3pfYZ6KpDssCfg2iNp8IuAmRVBcm4g55CNMFzHsJyxFTIdG/jHxSv6d8vXJZ/qgx
Wf1t+4J+xvuod0gJO/44KYQ9szwkIqulavG3QYWbrBe24kY/g1U8zM4RxdAqQFMRDakyXpu3jgDH
bXqs+2Y7LVCbeKp3DWixQ3M+dfoTFc+syZCQl3oeqL24ygnI5EOyXpV6nUY+Leg3PmqQ9MVNrndJ
1HcuC6WsTc0OrPdMR8H6IyOKCs6qclkb7dPJmT0SFwyeKrmZQPJXDphlLddywGyvGy8j9GLAdZUj
KkPpJJ12VLT90u7r63h2ui+hW3yML65zE5BoOCcTobfc6B+Iwpm9gQFvvQar1lzMSHN6auz4WtTl
yVQA8NTHRLLM3plx/9SxYJI8+lX9omLQzIQRAQ2OxijEA7NYzayMiSdAMNcgpowLvDxHpenUyFpT
SKOx8YJCkorVpnuOCo2Mq72/ZVSAD170nn4w2t7Z+RvIEMj7HiKsSkS/H2P5xfh3KL4UIX/iHs5H
Nq+9SXqSAkw7U2QCo3u9OZ+kHaSWztP4xw5LeUHTzplMauLEp1V1RUgeDhiMf5md8GfwANHM0Lbw
6vyccpj1z86uLDKNYIJa0vMvP3fTqyyq381E/DIHnun6yLm45f1ZSue8+Q/BWdRVEDnJ8lR4Z4CW
5Ou9wOw4F0CsHrxLx7W+Vx+DXflmsEZJgoBW+WJisal/41lBFKGw2em2sNBRxsO+cWegBlZLIhiO
GzixSPu4nGK9qksjCJCzGM8nI2UwW2ikGq2kXa6N5uBQLywNSRoiMh3GjOQoNn4qEgveXrUUqk2j
Gf+We4ECpceoBwBgf+Red0qJafo4U2URFzFUh2vM11QNL2xExy925fSd3419y+x52Z0rN8xItBmW
sHCy+D32y0e90VqYkgiIuJRZWajHXiR2/TT4UdCvwo2R8Bqcf92YGzuiGBM1tB2QcEoKuaAPFrF4
5O5GLYLtoNp911zoWAdHrKwqekv/7G7o23gNKwkDiTD0URcO6JGOXVtguqkq2mmXkVN0L+2QiqKM
3qV+gB6wg0kpWJC583oWJhYLNohNFggLk2Y0qcHy/m6hUUc4kC0txecOcSoUb2Him2pD1wyLKk7L
ksNQ5TglIJs6+U2yrwyrB9damU85Mee6e4bB4s3LOEz0tmQ5yvxBQ2qZz8nIXm9Yp1jlLyczUdQJ
Aj6mFKYG5Dhka1oj4ET5bKjYSfIzy77kEAGkUF0mUZOTwFD/eL5vWFZ2vFjTuhnYbeKtCxpB5XnT
iCKycZzey0cW+9kn61grqcaQFvHUuFIuOc0aUWRdHeqwR0ilI/O8wiVEqol4RqKDw1rl3vZ+SAFp
mZp6OP+5y97cbBO+sbEglAQaYeFWGs0DmpjGyaj8Os1RAllsLUxIj+SVQQFLIt5RrCma1FMyoO0+
I3Knkg8mGFoK0pQFZOhc0jcxHGFI5M+FWdsyD3PHXdRt10WkQef98RUTiD/OOEKVFtiB+fjywQjL
EEsph+TRMOMIoIDfAaNQtCECs0FRgGypM+8yaQj1ugOkvPWjfyM3leP5kKbZPhTe0YfhHln63JgH
hvkikwa2ySmxO0rlIxFq11kNTHKkEDzX4W7d44c8Rhv4mhS0GyDWRZZLv/41L/sZ5La65lDQYfjd
6m3TQeqpufu8Bl8FeWRGsd4nFoIm3X4OIIjX5G2J3O9sufADDLkfsQxJ/26j/aX+hXO7miUhD8Mq
CaEKFFPpySHfU6HD3KT1Gnrht1gyeIBocGu+Y1aQBWsLkEhIXu7ncYaH/veadZzgJawHPUmNH1Qh
e/OnSH0OFvqL5b6BLrI4DH6SNU28j+aiRgoIF7mIlBwH0uilIvYOHPMhz5am44QlZ+OlL2U4cccm
xpevP11ijFFMYPdPWi8AfjVOXBuZ4+ro0dlazPmQGEAmpJgxKT7+SZBJmlRl4FGp4sC4RP/f0TZ9
SLzj2cLO25WnHhGK9d24DUnmeImv2egjHXPFBowQcxpOKFxza14x6KC5oVQ+kqup8iJlTVwz6RdT
MSDPKJoAqakmVK7GMgXYwkjuux+QGHIuncCcectXYvPBUe+VUYBPY9BIYIqXbLkQ1fmF7pGjHFFv
juB9JLdcyJ5t0Vbsz5ffbhipzTkboWSPhHanzdoqI9O5x4AW77pJNB5cAJ7Bd3pU0ovMdTfOWcSg
VVbJEvq670hMpONm0gXXcSguKzgs/7vpbFQVGmAZqZqwYKbXtzwvDdy6tnjKtK/7hAFsALT639+8
iFzMnaV+Jk8smgXhKC6HkI12OdtE17aKodggWwALRon0YFoMro2y5+lQa241Er7gT2scss6U+vJy
lQs0KIv8M/6ZFoWh1877KClsUmQtTAob8+3uxthlBA9kEtsIzKlWMnTt5FcRcXUQS7QNjvGZ7Ng1
Bpw7a/B1AmNSJM2FiIDTtaKXiQO9GMjSesNbC6RMvq/dLCZuyI26jM761W7M/7k3x3AmhvHHmJ7u
77Hq5ODVAZkcHrma8eIVVEXb/vBpIENS1oxMiindfQyGFcetZDVyLBlwUGdJ/0WMXOPUF3VUaxXm
5rmrbamyJNm2V4g0UtqyVcES3eFGVU9WchIz+lX3UcsQimRi1PaOqdxfhYrTkcwsrJOEszkYfsyY
r7rTTI40ItFNDF7gTKUWbofkS+jjCN85Twxour/FT5aidYj6l5rnWVPvNm4InwWuRSrOJ8UW8dp9
WG9sJ3RqtkcNmNs/rtjgmkVdibA5eEAwWHrH77FqELbejznLcNugfh8NMmEDI88qRQ4vXJMZ6+i1
wv7/ZTvp/zv/6/cDuQBX9uUh767B89es4Pfju/wkTcHj2HsMS+uPAqSau8+biHYUwGSRBKVe3SmO
ScNEyNWCuzXgamCdpgsA2y266i3m8DErVoo1ZmaFuijz1Y3W2f3FTAQDDuEV0DJlzW9/XSmZk0OJ
d23elnE2cXqpmAI0L7s7f/w5CwYsjtmGkJE4iB7r5xVH6xX1ZUM/B7zw9w2XdVo2GTmCPPVsib/G
Y1wPtKwM+OhJe4jQ3Q0yRpN82OMEyvtDvtEltHy6jwEvlFLGne5bQ2lsu571HOma5A76mLtMwxdh
FrrXKB2NX8bJC3duwub42/QZHPy0gLHkXwblJzKZ57G8SYhjRScJM6+CdB/z44NNjhc7RJ6f2+d1
Ij94QoMKTFqfaZKU0HcJ1ffgSnncTRBeCYL3pdugasi/sSZ/1Yi6Uk/bQVjRq3hUJ57cGLAsCd/4
yk4grpTSnGWir3ORxjRy65LUnS26I4QB6t6Cbqw9YrvN6Q5rEEMIjAqvJUVB2V0feoDNaSNDjiwq
5cnJUV+FLDkiMRDg3BtC86itHB/sZmFw5ENh02ds/4ReC7rnrXuYbMsH/X+1I5NZj9geYPdG+fTG
QO3XeN8K00MnrlKqJz6JNLFHJOl06QB4aIFxa948XB3OrneCPbgYGsde/tZSf/teJHEqthx9g9wU
GkNYzuUFfHRwB3eDreMhCRC9Dnv80u0pM2RAdNy1TmcbDdu4VGvLfOA1qwdUQshV9NS+k7F8qdog
MM7pLJUyiFQxAcNoC0kJHchlvMakF2zYd5RTUQQzpp9/DJ+dmBp8JZX9cn6H11EJ2y/HWtu5V73y
oHvrDKp2L4R5OdSgpufMhV2nOaqVRzDoJQ3InKMbzza9rVDnsaEAr4426nGyMtwbgRxgaXHc1x63
LEfen8tkIUCo++MMWoeMWYj6W72clgqrMvqm3ZPTztFYo4WUUYiiOTrOfAv9SyAw47NOhEbqKkfu
bKLBIMEL76+Yf7y3gQIAxHiuM/nT3AkHnxBx3uTA/+pWz4wAm+g2Wn+cUp1ACVwUjyibUr0R+kpc
iEQOFpfNmYwUdHaG0cmmUZTUCy4lLJc72RM5RajRjKd2UmX9cr/wLFieTwaJNml22Rt8dOBw/ccR
Z01GimNmuay2WMMVyFBy7HKpxIeIqowQK+E/Y/qTVYdyki6A2cgXQUSUIXq6f7W4y/HiibdUvl08
Xr0kiUcniXYRBw7zIulFf3FsVzCmXRsViYY+BDdT6FaajZuWM9jGXLz3ZEYl+Se3GX9hkioQs/st
3b4Ic2q1dn1OfGk6pmdiU95Rq1gppSqx+tLvdMqLqh/xtq0JF79dHulCbhsBc0P1hHgBhMK+UiJv
KyquL0w/+q0GS/DAauy/yYQ5wS1l5Gq3CVgbGGvf7Evo1NTV9t1tRwkDSSLpswC7OonwhNVxw7FS
NGWtbebDQKTuLtcXcBTGtmwL+qG3d9hHOEp92KXK23yp6MNy2fXIMz2RP5WzVdwNZ72Fj+NayhlG
MCVDGnInoa+1SOS1MrcgwrdAmsaqB2Ki3bIW4xItYEPcfc6cZRO1W9Gp5JHbeOgv7CmZr51srbpw
/qr5YsZvNYbivv8cPXv+lXw9YAj4nxJbS3WmMUH9sOEzUoY5rRF9a5+LZ30g8/IwisjZDYtYt2eg
2ycr8nrG55Sz3t0aWIFKic+5WKvqLBLN7FDgnX5lxc437Sc+z2ZQ5VMKxlMIYvGSp0ENAtI4Ygpk
QIp70ShRCEp01gKVXji0AAwq7cfaZ1009qhBxPQNlO/DrQvjrMItPoPo7TmPq5v5gpPf4ZVTfWTC
x3RyFsqCu4AefYxGzvCw2c5NwS7K1lHGokavhUeO6HEfLwR6HRNcCC6v9+57yHbcjRORgRfDJwDH
15FB5xkmg62QD2SNF1um+I7Ft8gMi+JETDaoumQ6GiO3X88WrbCleUl7iSLU8DOFoxMa5SOTUOG/
76/zbBFsc5/T95hmJgYw7A5Uriwsy3Q0FI4I+A9/WAC9Hfwe0DaRpdupv5tvd4pzR26PinE6ptlT
BEXa0+1kj9wFBxO3gYiD37iW6cMY94tHHqnC6RimpGXY8klT+xmzlwmx4VN/AjfoZ75dMiMrmQvZ
OJfzKitsclJzqGmjgKNCzg2HoGi08WeobsVMxQK52JXOWPhRBdywBVgGKeZUkyWrgSj2Np/qfIIi
ZMAOHhn8K5aLt2tJ4wwVBRiOUQI+prmBoa+qYctdAxupwEByy7Q9svGWMxxKlnk1qIugq2Gxn9zA
hq/ZH5MQd14CulvuvExYO9BG6GnjfdjbX0Ka9R5RaZYyfs9wulY1yZLeRaOQfkl/DFN2zU2siw0n
FJnru95YS7w/gg/wKbhiMZX4gDTv/Z3ZNFqcENbmzZ5BmbxbAdnrNn2noXsN27VR0KsJHIYBgtCE
ftW0j28Vz+cNburho6/+3Gi8AfhKXoJFpXzeDkWqmB6o3SohTJilWhrmh9kQTcSwfoEu8D48jRKn
jvktwl7BP8Bkxr1ZgS4dLO6uxP1Bl2+8UpnnOsC4LkG0IPg5YgfpVj86ChwRRcdpXESUjT3tT24q
2D1frjc8P8F4yPV562EymJAbxzMPGU+n46oYJUBolW8ACVvT8vLvk3sfqwopnMMiyW5+d5U2NNqp
CEIpWPGa8w4jnI0R9T+IwC1hzDbEf4iHuoRLYZ9iJM7M+VeptJecUSMtNIHFBWB6aBd5cF6aoVKV
VQGXMLQc7gLX8/WEgbzfCTIK3mHFCdwm9bUsLf2Z3rVPmQPvqVONubQ0d1Pe3y1AUg/LPPjVApw/
4vzylhXGv71/Pe8kNgkVr5kGLge5FYQVo7dNpiBQKOuiA+3EJG1sJiekziJc7CuBcdDA2iKHlNH0
IvpQglHbsN/oo7sFw0aC2a4QF+CQAUzDx59mugR3FfmQzwY1TXHyYqzIqmaMM1EeWuxLV1fGl4dV
6N543+cYM4etWFCoCbaUwOE5oAn1prlRGAyHQeQXPAVOcJiBFsLjHrOGoZ2b3jZZC/CpxdURrWMu
jMdAIozRRjbt/o6t1xYZWQgBiRlpOMTLCUml2unLfmfGJd3FDIJoipiKSdT+djYDY6wQYMbBB2zP
7XIfHP9aNZQpCHr/TJkK/+cdzSO/fzf3mNeBOlQnv5ZrRSs3gd2gxPI+kMuXYy7KCNPUX/RLzcx8
RAWeVeds6j2EHhPs3eT9NvXw/MsjKrm6bJjVV/Xjnb97dC2E2hcE8cLVLmXK7+gtfjgZT+m1Xhcu
IDIXTjrdZA0FcyDZvnK1JqNwbQgSso+rOh0VJbIvHBkcSsOduT0CVBJ+eb/aUEd0f2fRv/mxteBR
vh/fSLriiucDFsuAHPj8Q1oOJFX4dyyJq2NVRKaIDBkCIS2AFrlG6FGfuZy9suWTqe+pCrCUmzYD
TTjQon5L67a94NFc+hcE40acWyXPrB+fHRHNcZN/lCkBevwv8+55O6aHU7DuGZ0wDWBEh2kY8lZi
q58esxDa+KQseZqTwgSlBlikQAAR4rJCQLVwgstnDMS3cL8xhXYXkiVR/ewYPC5KyiOVFPAMqCrU
y88GR4R+D7beAGBZirhfvWnXcqqIQgErKhQ12cTI0GQjq6vgUuvrjsHxj3RP0UMGAnJC2RoE+YsJ
XkJqQCLdh+dRWX2Q5lN6fpIUYAC6MS1Ul0DBvlYPf2gZ9t62lllyoIt4HsUuKV0E5Dx8W9H1vWQ6
gqv2Uvw02Ckk6AtPjvqds65eB5/fcAPQYS7fAtaC3trhnVPFPjL9C2hkdi7oE8VyQx94EUfLFLYA
2HK5g/qlau1URrepl+kQAUQYtHTXavhk94/MsS/zjzAaVjBEe81Ne6BAmW/phiLqi8vOP8372obg
1klX/6r36/PVrqOZQ8EWspVYHhRvUXIfXffTz2di1IoMsd64vbUTaQVxZ+laHBe6sSa88pC6e2Rq
hxmmd7Ov/fsgK3bFnaGtgUeCaYEphsVHiKLumtq7iFo3hqYSXMUv3ZWUhUZ+VN2h5Q1wuZaVRCRI
gjt7nLwLq7PxqmshrgiUMzHfOJe0cbHMomqdwnHpzJvndV69BDk1L02i5oz0anwgbPYxA3SUWg2f
5Yrw/CtoX8DhdMtkTbtU/8aJhNXC1Q1ZnU8k7k7HmMEGNH74cwCoCCfF6NKcYaIEad9sPNk3/g8+
tcJTqRH568dyPEyaKuMus/St4nBwbDD9v3jJSwt7Yz4vuc2wKeIMqz/Wmvj0LdIqGrj6TaJOk32I
D2P4ASonDqlrd6qnWoaMLS1CHnwI3VjmSTpTNd095WKm4ZfznShABzr3IGPzDNhjGZnX1m3SAx4e
gaSNxBf5kfh+bf9g+0zZioshMxxPJKVAPsXLHEqqjDx3rE5fOcwSBE0eX9sGG0MaTfgM5FmZUaxI
F5e+YetnjLjdlBHnvyUr2sVDfY4B3f0mim0tXcGxS22P6bBkVppcEvLozJX1A0afjQc/LAV09odO
Mx+mvFGs1f28zJhGCuJp3hzKrZMTR7X3WJ4tcnLVO7VuV/3gQMVlGuhUnXHbmlCYL+OR8Aft0R6j
hGLUUO+qgWgv+JmtZJHhLETj0Q4EQXhJyrxMzeJ5Cao6hvGmS/+Bu4T+alUmW1H9OcElmX/uljMu
U/Ygz38OhAgG6qJqMqlnl/Y9bwxYQKndFiPpR/cUjN7KThUrckkyqx8zWaPSiHOl5v6xXqfOIpx6
PQClGrZ8r4nxTWeUS0Fa8KuheFeVOwnzv+RiP9RN1fJmIG0CzCP9uQuA1m599dZ4AFknV9VeYHDx
Pu+FBBNdDM/FuZhjQpjGTjibq+3/iv59uW8RT9F9pIxRRwIsUXAqrKixoP8C6I1Tu0KrGiQHOn5k
gZooUCGS23fFNAP/bg6v6lZ4o97Zl3bHOPITBZWdpB5L7cIwbq4yFvWufKSdD+C6NSnO9E9q9zY5
4qD6yqx09qCIKs88XchuExmFv2ov9etMx21Xl4pBw8Tc2u0dQv0KcEpedWh3tgtaBeDcG9NJdcAj
Tuh6EiWS4bZP6xIILwjhA+BeS8rf9B4SxUeb7HJaiYy5iS9AYaW1O1Qy1G7OwkNcAwiwvl+kOSI4
jhI/chXLVPWC6WeAvbUc3qLQJ2bjX6B+Ds3IOSAYoMOaQ4H+xQWDeNKbiZ+g/nT23K+j0A7+bHmA
S77OTzsObUFkl2uWp19mdGsIEnDnqiclnuMfJtb4LuwYkoM2nektGp68EsKirKbrqusM5HAE00YC
Nsz6XLjqOfndVzD9hq1nidEF4nXLRPrAqfq1c25nzP3FmOtkUCUZbZAIc6lnMGSslfdKFPxvMozC
WeIoDOCtlstBaYDhMRht8rPH9L9mdKXXQQF5JGH3kbTMp7v5nMVafwDIDvIv4Rp7yHoCA41Sy2rz
snQr1sqyzvHa/LDBHR7HyubmNZMu1G8BhxinQw+EUwTkCR5YBeKxhF7sYpt6STBE/LVNkhPIY1Gu
U2zoLJhDq1drHLLjZV8Bel1tUPrUUBcfxouVZ3UraLTAOtx3HpF81+SNIInmuEZxP6oW/XRCfn5j
UwAhZmg1VbDxb3y7FLWQ9ilsmJ88wCbgE0YvGWg4QNtkBGkikg728hc7kW5d8b2xku9ppWjkkJ7U
xh4G2MU1GLOo5JxG3uR52a5h/NVY0YfLHxDJ7pAItle4TlgBNjiqxEoE+LRq06zqE9VhTvVn50mm
FJpzjMrSun/McjSSwMq4mKEMQh1MpjDpUski7rAeE3pVn5qYPIlVvu8KpRtL0CypkVew+Wbxr524
3U+nWmZUx3tUgljKns/zTTp2QapCDDmTHGxS2250d/Y72UBEJoSOELBvwdqKkw1gzuQI95SGejrU
r3nQ0+sPUJ3qYOR1fzouTXIQNu5LeA+8QTJ7bb1vzS5Qymgo17rNf8rpv/toRunXvV8gElUe/CNR
YD13WgdvNt3mjOd+29CfjNZFS+cojjQ23hVDl0sYS4OmlAMAPJm5cB+vnEsOTi2QZNjC43Qmptpx
0zs5oZb45ENY/KqbFoKwBnvONHF6XXolZNCJRxa51nprZ03GoDdsukYTFqCuK2AudgVjyzFH6O7Q
Bi4l2k+6vLDlBryVv544SuJrd/XFkvmhR5RzMY2s4PSeyEP8Oy/gzVS54po6fAstbZhkeus+PZ16
nL4wFP2TUQ2Va/rdwpt0jE61nSI5SJ7cT7LBY5xHv50BAQsBtEuqi7TvWOyHG0NtwrdirmHz4w/C
8iHzkYiEGR2zuCutntSNF41e53kNuOqJjd3B1pdwE8qDAGZyoAO2Wd5TumEN3TWDIhmxnXwY590/
/rMz6DY6rPhG7esXP5CkTnHKSxXeOXer3YxGu/uLf3v5DsNe/2ljrbgAwKd/ODx4fDJcHzQQmobW
5EHosb/UnQByZWCH2dGBcBuUeJjR8CNsML/iI2Zj/TZM5jDb+ovMtfXftoQPHaowqjN6CzYYV+Ja
5DY/Nc0553a6Iqv69Nu3pn0Q2Yj93ZRSmcpLPOSNlwAFqjS7lwy2Bf1iWj5GInLhHaJ3lSN+M36n
EzsjR4F3nkv46yXHdLa6aElcG8MjiVlA/uXxu7vwr07jbPcR6MbpKw5TzFZxfLIbfjQ39UFsneqt
DORncc4N0OYnsypFQazsFbkztXeCGMa5WtucSmJ2T83jWh1eb4MgnlBOxgP1NJtdMpyZDFRwiq9l
fRd4VTM8NTOAbBhFlFkCHqxvMqGiGVfxpLDG8IZXfzLz85ybPHGnEZH0pLJE6WVoHMjI1sOZ7YHQ
gMpwmVCGdt26O+P0bt6n664b/vL+qgIKURZSACJCLXgtHfytx5KoWcSfH1s3ajletvqmIOVKTvZ2
fpzuouxfDrVPayqBBQeAMlY1FTY24uOFqfr0k9IUb4KwopGo1X2QQNSnPsGHQX909aSSDrrYHytl
aVj0Cy/lrOeKumqPug1RKeYO6NISMQesnW+FxA/DIy6Om4/YH2qB3q64b4vdoF76aZNIY5Y04m2G
+MmFfldJyOwGymKBDR5xmrayZ8MxPhupSNupL54uGeTkTdMhFoj0sDv3RjHbBfQdXLZncr06piaw
SNrG2HZpw085lz3Pm6ccvelb/YtgC3YpsbuipbvBFF7n+iVnK1OJ8yGhgHcVQP7Y5LHUmxgV1RCo
0E45RGNyZ/Nj66LleN/ynlnzkbpKfOtrSH5oLAnDk5D3I4sunsjggcglmVsEwhlMOdOC5KUr4M82
Fo/LASbF4t6HL0d7EcWBHEcTpsEFK7nVmcuHElnQ2lhXn0EZCiG8BeYKjPb6hpESW4hAQVzx0gk6
bCUo5VZ/F4+JSqHTdyLwEil3J/e4nj0gpdzur02eLvwAbkoF7DVYb+K1KRgx1VOonbzgELZkxOWj
yAsC6ToTJUW3R7BsJHd3ZIZuseuTqEee83v652aRalsNiNkMtBjgMQB9KGOeY2NaT5ou0Hygmgvf
MPzUQg0p6sFUFqMxkO8+pO/Z6sxQO1CQxeKztsmxms0N22xfCCdmddwu1EodEdGsJB93PZ46Ib92
9QZn2Zn2n3QcpD7VCio2R8pubMoL0+KL3XGKW+H71FaiFcPe/ns5lw+f0L9eCcNQH4lZWUuVm5Co
AAqwoftZSC8fkTVY1CsjMPJJ/XHYoyO0hZhqshq29S27cLYggTmpbRFaJdjcZ0uwXrLyKy4Adryb
sJDBfdyQfgxnsvLWHV+zS4MerEFgWbPdRRS6YYFBjIaSW5VIfxJow7bJdFQarn6gChrt/+ivcl38
+azC/tPUv+GkKwnr6rcmOUgZe+JyLRSC/9VptJbkZcoAh63Q1NJQPQ0LNniGSGrxupDEdzMq1GhV
j04yWUptrx2AIxLa4M/d/LvuZ+YO1ZMViTQXczKtUoYjAu5aSY/08+A0b0FSQj5Qj90EFCx6jEWf
9PAq49qH8CPVxj7FIxsk9WwrJedr9tvgIWRs6wQ2Mn0KLRif74Ndl53ZVwQM6lR/QRrGrS3PTUE7
cf7YCPlEmOUBJhlHl2sF8KabZtHo+/Hulu+WbDuTpJN62f4wmBun2l3VFOjex61wmgOmihBkrz9j
fIZ5Sspr/Ka+O/Lix/LrcJyA+PORO8h7CIId3kLed0NFv35+n73Wi+bG6O/XIQYhkz0xmGPnondf
Fiq/wdJjJwTt8oej9QtgMGmZ6sxPtRq6tXtLmWcgNZDz//8tYKc3vS7kdXbsbHaWKEPA++OYjOYE
N9XsDAt+PyVQZA49YV7SfJU1qqOsZQygsCygOvGb60m5YTMJ4ksdCU6ajNBvnSYE/8+fkeYPhJi2
hCd50xkCZxGlmel3/3kh2dK2LqXaImJiUJaWdZUzNOdxaxCj3oaF3gP/msbfHRJTyY/QpYiByF13
cmk8vuuRIH293OXAAEIyYmrzdv/CDM4yX+NQZ/qpFFNQcHjoYlxfBXplPNvZeraGrw20/q2twFRi
OFdlxtucPYDSNP4psKzgOi/bq5vJoeL/6LKOjJa898D8o8bnMMRV2ZHi3ktsDVI3Pi0GDaFPPb9I
9BYN1cH4fTDPhDvVhvDma+e02KuZxPqOUwDRekFO4rqgT6OWhX9dq4omkiC+uIr4yZ74orBCzMSm
i9/z1L4gk0aZSlPo3xi/FRG71NUfAqYhIIPqDTtFo+xOQVHXi3M54yyFQ25wb4hO3lUIbdrFxkjp
eNfzKoU/dqrSY7WEz6Vrb858xih9Oxj8Tu98ZTxFqdLFjUoc5J22kQ1uajL7kmcBb7JFbwX08L+2
Au0yruPO911wNRE+tH2Ggm9RKYDATeFipCMMhh3aJrH4APRJW2QXKlT7a2Gjyfw06pRIMzMlb9yE
heprlWOwxoh4DRIXXIy3aFTUQ/UtADAFXM/3mo8pMhxAgl8b4QoZL+Uww1HIEPQgQfT03/6fFtay
mJWzDNPni/MJzjN8o74bBNS1olT33LS1nw83oitnY2m8NyQ+FBp7OtBz+I74JZByY/e9aQDDWq31
skec6nxI8DkEpykN0U63SAofrG/wwKq1iFfajHAm0EYx93rice8TlW8F1HFgY7T0wgfbBay1bgcy
xBl1QO5C+7/z52k3dsJhfvcuNm6he7rcnQIKPBA6Kmcy3U4wuGdGIkZJqB6ooAy7Jm00xhDlBqDQ
gSMPrOvNa4teUtrcbS1WKQrQyR02O1/Qz9cB8b0oxGv/vu6TOiNuyPT3ADzeQJfxYPxMR42durEQ
dCLLDnFLwvHTUwbmCKMFYFdDWqh1z/nc7awrtZ+YJnxJu3MqTpGvjRegL2VeLG0phH2fRloBlX02
P/gOvAHTmXTazSkqsMdUTZNJ/cmFE/kxzm+KhRDuFDG12L3f7BbNvHFyk5soc/y6KrDPN5+fMJLm
o5W+uQfKT3uvA6XJX4VdTWXfPA9FkW69WJGzAaKXV27vqN4jFGJO0Ej8CXzKfvTCAZTJXAYT+L2x
isb5Wfz20E3SNKDEUrYFviOEeljUhlLd82CDfnJYNEdNvR+LcsRA5tP42In5IvJ/G0jMyLhiGqVd
2c5QFwmySP87YO8WLuEji2SGIG7Fz8iWRcCjApAbrUAH8BJlWK+EOqniX1g1sVp0AlhD57re7MsI
My7TIIEg+v00g6i/bl/7VGYy7LNrelThiqU3PbR0LtRtr+kd91ceIu+4MdxAm2jTB01jLxv6stoQ
KOQdNqTkHh5KtPcP68AVo5avltPApkOb9Iaef5z8x+dTTHdjhf7xGjFtjF9KdDXO/BqXucVcIRk6
Y8mHeEjaB00J01vEYd86+HuIEcO6zkXdXXLjtEOzMhgT4qPG9ixh7SJu9A+FGwTE26mzf0OleSYh
h/m5iwyza70JQUCx5e6yc6AanG0IDS5xS8/vnsvhnhgADGg8pRHaiQ1aGkOQu/tob3vJvHO14yyE
7mnPNeRHDC0zGr3eyQL1stQVray+HO3WtU5MOKsi5O/A4pGXsOTkLqWOSTbARVUFnYn3bOw1W9rp
2niqPv/s0C39a30GEvNDp6XvTDHRG9H1ID0DAaeUNexQ0PVoPRe2wKUDj5tWHXDgF3paMrATKQ1B
n9pl2QA+GTrO98eT5rdE+IunIqXJRJbCYRzJ5W1Lo4zJ7JPiabo0UhkrIdj0KNYOt1RKgeto0dfr
Iwrn9tTTNmwTGflH7ZJ3E0rw3N8gLoGFGqcCtJuTPp2J/9GYqlHcDGEQulqn1khahHBc7Qsv7mDX
AQQsUnEuYJozeUYCENyuKtMYMgKartBgZ8OkDsHSOJDB+H6sb/iW5Onkg1g7DYW9jBy6NCSf+6Hj
Z+vagPMzxnJCwjN+2ZN/SWrverTbg54u4LWnrXAKZaolVUcntKmoTgQvz/74ToRnrGMnlJPFZHVb
tA8+IKy53RcN1MJ5E0/QKeY+xd1BLdV/n7uNgLulQ7cXeELdbMaFBGYNWxoIEHMf7y3fcHS1JDYc
Qwl+o6YA2XMYKnlwfKKjkFudPwJ8eEo9oev9duMNwAHtY1b7DW52eHYnpamk99wqWAcmkCu5vu2v
+RFkDxCViWWD9vS/YztramlmXTJvNSC6QdSaMDSFZPFgd2tRMS32dQ97W+eZuN6+x30wGtrWYPrc
Mlwde7zXUny7nxg/cXCEmDKp/RUUTI0IRUi7uja1kTDNYK0AIZcp6o9XVujwdMgsp2ZJZ4gs6j5c
EOD3YhZ/B7bgaTjAF2A0iSV2K/04lxLUWzIbCHwer2eJspQ9HoWW8QTDEjS9pPz3cfob0fF1sCMp
Runsp/JaQPNxPRMSTwrngAh9X1zf7qxHuVM/+B+QMwptGDpdzxqaDjVNLRYLUFomW/2Id+YvywVQ
GJuxH5hw/GKPVqdLPg+CyjkE5xMNd0SeL/0n9nC80J9A5bJ5Dl2gT5P46evujb2bvy+Q5QiMwIQB
Xra262V3/nVtZjagW5FfZi21CHjLpbvi9IARgpG1QdFyPCEq2Tn5hWoOy3jzslHXeG/uYiA50hqT
Iz1P0f1FWq58cjuaxEiu7if9ITvyNB6Sz/WFgCPB3/NrIXD4vQWNTSbpZLwsBlUK1nhRmGexcKw7
E34uJmIn6tRaXY6JE7qjdUy7rUeV6vKJULQOJGdLVC8bsI5/eFbv3zbkd5zhKlT9MFvfvtxunHAi
1HNEDxpA4TTjZojONwDQuyMipYdRZDL7sbLw5vYUaYyx/c7AM9LjuezUU1ofRoeMKrSB90p6rO8m
zR/wm6TnLzNQ4/UHxtIfXECynLx5Pl4gDCnHA/zFV0GTBVSFhbcH39jO9TQJ2AuiKJiCiexCxg8J
pfJ9AHJlTNOO4M962TdBErUbAMFJ5RF0q+RJqz9BYTZ3tp9MbD6giCavHUxpyJzJ61gsVP4jbyCj
6+kchy6iKdKvcI+6H3n5o/mEq3mNnZ0/P+gnCRJuQVlhIcP3uIiy37zfaEciPoJQwSIEmYTwiUml
p7zougABIqz/EvD5EtO7NO+1eMs9ddzAOuGCJEXgIojhxKl/qtdY/4tdFuEF6cOLc+feh1yOwclq
fEs6hxu8z3R6fnusrZ2qF2C0uqbWVE0IeflAcn20ycyxwJ05O2ZUbM+azSsDezVsnFPWUColMRus
MJiY0DR7A4ms5iUlmTDh31lCgzy+vTvmA528ICFU3bSbex/nv59wOpUSXyWuRmyWnCoWj0iv0KZL
BonDbsKR8Od3h17vVSNbYrNDDCRWXJYAD32Q/WDTMmCZpZOlNDlusDIAKoG3BbvmakIfUU5L00d5
d5fKra1U/XdQaWOa0CJo7Va50xo0v0AC2h6LKvSH12uzLX2zaZENd6neYDQmet7mfNtxFUZzsczT
CAVbgmO7t7PZj43Y5LpmLdUY722J/NcW8LF2Cm3zWf88mbaNY7VqPNN+PRXNunOKKMnRCPE1CYVs
AviDURFFPlC8Nfyg07gmNen83BdJQ3os5xZmMmC4eRuvBTUwLqilBw+ejtxXznw+lpv33Zh8FeDg
+jsmRAqZxB0zElQMNwKeo+s08KlMnH6rL12fqWTIJW+zjI4keWtXKkvRSZ7c5W5E486atAURA5Jb
8pL5QY2QF42mJCwm1co2JvfN5h/ypjBuvPaKbPXWmuJi7o9txlF7dWtom6dO/xhTCmuE3DGg2II9
UNPhvxQYCFJWAdI20cVFEV2q+zWBIrZqmGfsRsqTujB5LDHohg5mW4SNEkM9TakE3+m6FRlA08F/
apg/u8c7E++uBRsYa0J8ap6n+b5aRu0I1MPomnfbWVr5etL1oB4a6pGz3rhxhQ4oFS4eN4cA4+g2
730I3PU59hLOD/qto3e+1IAM4fFMeGiGkPtR8iKQ6xpUeiOIzVP3zpEm7K0KJwkz8whob0CKb2ab
NYfs3lT8X4IUQRrUPBTrZrjee2DFo1dQqHif7lrbkxCAoxV8zs3YLNaKUX04qFhAGsPUpYnVNZqC
uUa1ZXR9xHvnURBRp8AnNEZWjwTo+sjFLpAN0T06jL4RkuFN1qTT/a2/nQ/NPGZmQXDBPRxJ5hW6
foHBt+SA3FXoMhfcUFTaCecb6r5GcMzwhnj5R7EPwJGBWTOKEsiNqGU85ghiJQmfZAC4NnSJKX91
VjtBqZR5qnH5jEjxVZqe0Ns8Bi8w5RdbR5zmcv+vq2I/2d1lKZ22Vcd3tgbPqu6gqoSMf76FERZd
Cq1K6RtHGTeCVk1+Z0uMRM+OBjkvE5wvpYowMlcUmExn/Xhdi2H6veukZTcC3YtP91rjmYXiaeQx
SwFRNpywBmaaM7OY6zMgKwXwhUxnHezYjE7Vb3Yin7SlQX9soqhkGF/dUw1ED/1eK5MlhkmCW9Wk
907G5WuI6SJ6Y8sRinZmhLtStmFARpwggcW1qpQDxh5xcSKUK8/120kSvwgkcJ11kasuzNBew+SN
Ire4TxOH6/IKWAssb9wgZwgoXTxRNGMUtKfcG5XkYHalogsmehgSPf+tYhbSq9kQQxsgh7zY/TSC
B0EpxI5zkjBZvPLeYOrDSrQKLES32Qydx85loVn1kPC5d7FymjasJ9ZCWkVzbT5VFnwKbN62ChZE
q88+Rl4mKg5rOBnlO/leZ4HYUqdO9+C+SM0iZZOFxmOnCvjb9mInEFpXuaniwLqOCqrPEaUKMmM6
NUgQsrNaCF0Hs4DuWuW5S+D+I2QTPjXN6Pp+mYgOuXAhwiBQQBpEelfZJx0RsjCHXVh/7fd78b85
pWZ7+4vrYCGMm5GQRd9y3FBzFUXZ1IRcRgqC3Vj1uNP0e/l+l1tw6JvvI3ZJDZlT6g9/6ASaUgYn
ZF8Vrwv9VvhBxLExUx+vfyl1hg8/wD4F4lMXibw2s5hIx/hnXxreqHtku5vbBvV2vgNSFMoMOsr1
5DlMV5Y8BQL5dL0NJxz/HMJereXT9PJxnisUzMBUbZjhAiUpAzfXjguNdavkvj/QrA+v4fx5+Nyx
wcm82Mtb5SYvmbaf2vZTb1qziQLqSJt8XlI7askj46JyClWoaY1EcqQ3HysUhsFLVKTlzKcRKkOQ
3J60zgYx8C2Cu78fy0VFvndh7GlKhAA4lDjWMLyADX4oR6OzJziOlIgpipXO6U4YJmjyZsfS3Gf9
ABg1xSU1ak/DdIusMTPKP+fxlxovT1yMTmSzoYD6sfSqE5b4LfmfuOVFfR6fGiR1gKh2TDhbqYyp
SCPKAkigEYwHlFFp+Sy0cCuf83+d+MVvZBFHoyqZLzG73QEodJiYD1GLO+dHH0Fsn+b8eUPxBX/a
r93kyHuM1Nwshi9e3rE1KmsQBZJ5mVxlAncbTEuJZOqk1SCne3NcPpAQmeuHK78KibhYa5KqvLyJ
eXgH/+dmSdbe1yOtl0pEhOUvAj+ayA88CNnL+raQdYxdVsdHVhN/wPkzYdgJGHT4vlHog03bek6R
EIT4eGs9k+iQbkN8M4+6T55Tlx4aR/zQlnYgX+CuFfBhhP+2ilWP1/JRU2IZ8kcQYoo0hK+tzZjD
JRHDqBDs28/uK92AGNER5G7kHSa+cDXbwHUXEVNUE5p5jiPzOzwnupFVIZ3CCMm852G7OeU8R0r4
ZYxoLTR0bCuFrUHqLJhtFQSsTF6MiDyKDotwegUwBxmQkkB67W6FMk7XdzjTyT9GGdhkPM3FKLB9
ELalHNyIw3nJf3/w1/Tp/F/ED4/chCpGM/3wRIz7L3RIPZDC0J9RYQ2BS3THXAN/368Lp0fHK7LC
/3MxiicpM7LKBy4wOrnV6dqcjVGwgyu3qQvIBuOO3r5trQTu9i9C+I3dyFcP6DlDbANZO/jeAIpS
3Hded1uaBhuA9/Fn9eku8OQOWTT4+WpwXfcKf6bEp1rECt3uXGHkkC+iPA3t6sEBx8Sz3sfgLnIU
KnRLgsKuvzxRIn6cyZNt2BAkmEFsJ5E8SsYcmriwY7+uxLIqzx1df4q0b7LkIiKG1lNwzNjsbsjg
nqz1Z/fvGRrqRMPUagIGKNGgRE4giNA22hEb5mKwF/OsQFfQFNF/r1CauOIME5oI6gi9KfaKP3bR
L/Fz0caHHO2Rwyk2Yy2vcmuF1isBzMLPTCTvtFe95aAmhlNj589S8qitSwLZfx7GCnTHuJg2znwI
fiuReAa1f6C+cPoY4cjchdiTyzMMzrxYLN+RI6UD47z+R7qMdczSDCGBKLvEYhxtyyGysgZc9uXR
KzjKWjtuuyVtGzIGCZQoYaM1xn1v9fg+JYWIDH6XunFfI6C07d14Y599EroM0ZxXw0nJVw70Ec6K
h1MaSTMPjm3y3M6PmI/+rSNylw/AN2AmuvWT0Q4cImkfLsaBD36LQTZnoOAg5K74Wqh4uZLX4EPT
pSKEYkXMpHQiq7wnRcGLUMuz6QMc/BpWxmXQq59bv5TkPZroYLDLlh5Nf3iPUf7rMWvdE2q0Uxtc
JAvVftHPA/1ilfCPK+Z3n1oEZMO88RYUM5LrTqCS9ZZ/UnPz1x+xRIxWhLWmXlRicrCNB0hmmtws
ZfWh519KiDKT7/XD/To2np7UuOmxtSzMJtvfph2J8lZ2Ypiwo2nwVSRVFdaSIMPSCDI44VFmQRVn
S29mkGEUzaIhyFGQqEnDxJBAVDThRowMtgAmM3BPOw0vXru6vttjN9qvjaNfc0VUnIOLPDJw1kvg
bMQtgJbnmbIzAMU8xKXAXJ//UHG68uoxTkwzO/1aEYfyr+462upjxU55q4jZJF8PevIo2yUFkb3s
QFY9TnevzR59p+7jZ75PEcXoWw3C+6/nLQH4E0KDQGmX93/Idkj+MaM2iBJyuUoJlL2934ldeONu
pwe0Nw2tcwrED/SOIwbatx5Q2iJJhZRcaZQ9Sc1stSMNaVIaAoEGIIcz9aChnhDbGlRsYvWb1KZt
ErouVHj/B6p/CPWZLbfNjq42TPI/ineW8X8JuYsb/HwRa/+zohWBxd8n76BRE0qbWGBe+SmdPEGY
Cz02R9ka+ERLQUI7F7LzguZzeSItNeecY980K9ghnmFIH9r6vnK+NufqIY+jRFwZf1lXjI2HltRP
qMienGV4GHVCT9jZhwtyo1DBQrMYhAQouCnKJjWKAtEqircdGBVHH56xtZDFqcJwNheWwzoFNo55
DA2NQtlVBlxPqDyRTVsEWU+0iV/BGeHg4z0IQoxyayPKvWCJHXcKX+8TPi8fVOfi/etnYvx05t5n
KhPpxYC4Sb1w745F3NABQxIlDZ3RXuZ5+HYeD7x0/3pMGlcfASZjV6rzhd9lMMmfVmGzf0Z+3B3T
KsV8L3vUo9wz7q0n4/+IBi2cSbJ/V8ER70sLQra8R8/jKS66+xidLZibzFPp8UIb2tzoUdja0CCq
i7wIzMjLfz7s5sWBcBAHh4crijypaSnUv/cdYF81mvXIXplgi9JcUaoHRG6Qn/cXNecZ5lZp0tDY
Akj7ADJKxcWL1vMDF5NpA+LevjYoMeis04Q2IDLfzoOnE1wRNAR1Eiyylsn3di7Qzw20gcpUgr/r
O8usQP/VAdHCf/PDtImuq13WWeBQba4nVBAByKmsICSQkib03Y1Rt5Hv0UB3ULgYUtsC0BwwDsXY
vRPA23yDFBpByrohStj9RMxJyogo/mGg4Dejp7RzRrnKlwcBxQpZYasGHsAqvmpwgDJwKKQvhlSK
cy/w9BJEUEdLPwudNe+qOx6VWBMsA+M09iJQ9Li1lO+3XrdER/UHtA18J3sJZDIeI3CO7yMuySIh
SzEhzUtrjBvi4nwFKi2RZZheevXHKouMzjQze3TxI5UvZBGtF5hNFFG/85jTIr699eqXANP7BshJ
BHnvGAJfBSKYG7JDK6JTvHrvu1AsCdX+O3Kj+VuxRAd2iAu4gP2v16agGAkN3IopR1nqRejZb7jJ
/umCfVcriWnfC7xomdvBApc9cJGtfRoTXvzHJfmEpOsCQLJjDcSjXy2CJOI9kefrkxD+Z/2gsNFU
D859pQzTzFFzR0fElI63is0JU3ehAvTnj9s5591wVXLp2XaM9awVu3duehfq17zy/3ebzqOa7agv
YkMBjHlYcCfctlyxAqo/9dzirCsH7cam/nU9iJ6tzEX9vrBxExV3e4J4jad8Er4Sb/HVUp1QzIsH
hTfMrTzvBHdAvS4/zNBN4joS5oiwAsgLIlDg+IAroV+0T//HmGgbyx1YrOsRXshbymQ3DRtvix83
7YKbj4KMABaiHL/SkucUDmRk0LIVi4RGSQWHNp0+tQqTTWR31MSXn7F+Qz5fveZ1swz5XuU/5Qdy
3xi3N8Y+8LiTRwRV9JCcggH6JBaTFgKa06ElKr7aQab3WJE1rTws0sBCPjWnnnVhchxQq1qkBApq
LeSnYXOGvTnejjoxqFnx0W/CdWQ1jqO3eOIn1PRnpqybAjM+UKOVFCt17PohDiyMV44pb0bpAN7K
7/pO0rD///PGykBFlbIA28/NlE4ul2iYyhVGhZaGsP47nyI4/23eomuZoVxZe8jqFGIUnkLEu5CW
0WUZ8hGAEIolgwzL+jzBv/NOYtk6Iq2CsnCXgheEnejreljjYgrbfb98qmIWcbORqsVnr5rGCLJD
wZD/tADaZk9YRgFyKViqpibNRgIaI5edBzBsYQ1MQZKR3dU8cdf1D0p/SJoRbND2yitybBYz90JR
QZf6R9BDtHgzxOefPKHvgLwULowoRsmhhnoo3xQf9muX614wpq8nCa3iuTcP/EQaE9nHVC3SHQyF
CsWgJ9HO3i09s0fH14YyzLORt9JpdOOT+S83zuy83CsH6taKllk4Gc9wFYaiw1yVXEq8wMQ25HDY
Abfs5Kp8l4P3+PyOXCcu0OJzIHdtVoRwZY5yGYxsYVCwVP1HQQMiFkdBqLcqw9YxnLAevLow2dnF
4K+hdaUpQz4RwvUSiBX/pwh85YX8w1ts2TB+/ncZoHt6W6Hw5S6EhqRWB+uqIY0oWXtEUadRIgNo
rQfjEQZFYDNL+V1yWy8mJnK789PEcU/mc1HFPWM/LiRxY4QU9HmTQzgm+wanrsyuTl2Fs6ucrfXM
VVit3j9iTPLFbC18rxOd37JPN2qnseVfXJaZJu6UYVEv49r/eyrPDNR+VTaUydwZdvUBCsS3+uqE
cAxFhswSlYQBVS8lLXmUy1A7sPxpYT+agXJIrjAbDPuU8rArY9+UNVyU08RpMWuHDCEcyrUCVWsj
YTbrnQn5nNRqPpAfA4IN4WY5xJnjMInr7s1jrCrrqU0put+dOZePQyZKHAh18X0OHCUTpUxtD8q1
bkWwjV7B9i6NDHg5ZTkxCNdM/bj7DPpd8vXnWIzhKAqtRhgSene9RBp/YjZ2mdztXvD6LhyJvOPJ
pT96KOMP4SfBjhZlKymCwqrTTbCIG7LqdQwU3ff6Euckf9cgNRFbfDsTOYzCXnTYZ+2w+uDQo9/u
ur6/26TISYfKI+fvU5UAGBMxDtLdQ/rNpkL5szBOqAobHMvf9D1+WuIOF66F9azu89rzgCxeYnDW
sQmybtdkwdUZ85008vdrXJrx5Yc0ijnfsOQs4aqpJFwi5XB89KfXNBOedDKRaYVm4NylGkEqCYJl
0hRpZY2z5mE2rea19j0PLFtCruB2e3ugPcUDywBxXXFTh0b+N80DmZyTaDMAAOR+PpzUGlG4aMpR
EFvp6rdmPJ58dM3NaxizKKRQWZ3rkAyknuBNkyX2MXacU/TIItrhD1ZmGAEUMCzOKy505zPAQ/tO
iDTIXVkPLPisyIvQnfFBI/Ebt5eVkxyrkR5hi8LoYgn0xWF+bthucVRkbeAak52qRShuzRBsuRJt
KiG56Ri8/32gFka7R9Wt8e54kOXdjvMTwysXo1TOfVI0HciLoJ212NMRSuX1Y1gDz3UIC3uFDz7w
gCjAKVP7aNfTydVll2g/B11fLk9XugMXfQPml/0z//Cy8GDMWvBQoxBmCVOK2KFb0MbLrqnMF/5c
YTLbjq91R5pD1wbnXmfa/jyzgrluPV3VMwIRCRlWDsOVFZZDJc4GrXacSC+UMDKFC/zAHLNdGF8X
I8zQZJ+WIYByZq0scZD+ViSZQhItI0aRLTYgP+MhZUObR5geuHuSRTji5/uqKjsR3XrJHaZJExIU
NypWhQ4weQjtzIxUDwsFAKC+Z/i4c+QZnG/wEAcROx8qYAdIOL6b/7+hHJmywUWvtCC1GzuuwarF
dzkfcB0OkpAvq8PfmIcDsMfOJot1hj1S2NjtI3A2vKmVPiB9Eb/QHpZcwnzGT4BfplBWVZ3+QWv1
yJx0Cgvt6rk46WPmV3+BR3jf2eZcHJ2s2mgK93fqHdHDRz38ufOk5jLSDj8rHPvzx8DshcOxj9/O
3Bx3QDRL1kTUFHl4ek3GR84ke4l1beA0pxB5IFeDVY2647s9h6gFR+WdU/EC4jMVW1ytG3ynZcVZ
TnEO+IB7AK2RJFCb9VNZ1ChfC+O68AwOMj5a46K1F1Xv8NmD/+BvkOC4F7ElEzMKnpS7EWKd2wt4
uWQQJ0Re+q1XRaF4hX6EPUyDLCCSpQrdqYPB/D+Lq2i0TGjdvcUKGidHYb986hpcDwONOo2UwVjQ
TkatId+b9Wsq6eWIMD+8KT8beJCRbzRZnCvJsZKaYohaJOJiVaTS+mw+XUMs1yHR8bPAohHHlhlO
irzshrmKyL0keQj1XFqWW3rKK/z4G9Cys53RO58JCAk9qX6dXfajMRSZkC91fHTSgIO0JCum8c37
SHeq7ARLd4jwg9+pn1qbtor2tZI4fahVmVv/FSqx3yxoPMFzqLEo4v0Re3qO/jZ37O3HM/qUHe0d
cwRrJ97LaU1bMBieLs9GNI2El/RRdCvnBGuxqI42nKcxr9Y69zEdaWCIuDKXyQOBEzP1bP2hhI7Z
IlDeDS821/AdXq2LD9E8gfjOznVuLLkVRFEj8FAD5chOCseoKbXzP9UPFkBNvf/0kRq0UEmXAt61
cHwuj7BR80vhTxoDHFNQzXOArUIx76498saxGoX7vFLIJCQP7ICCsXwGM8NHSHu1cfW7UYeed76J
9yzwCafI9rItYAZNMb5w8qQj9aBsi6Gy2sbGnsOb/Q+VUe1JABmVtpiGoJf8Zeq0I9KeTw7r+CGY
qF9ubFotsB+YpCo74RstsvR2hPv2BBO2gZ4RVhxe1Tr855+XpmnlnmD5Efd8Tx18Ht7qruhcggkg
Bfqg8627Pfn/shGLWqdAYov/z1TQPwjkCqobcYTakEPuPcJjPgWf6XqSWrIZiTNG50ACyrZZdWBQ
kQ38b6VHd/P9+0D30gIr7HHeH3BlzE4tWHw6M3UAFR9gdfGe/752mw5SCfDF59uS19b0GzQTk+/0
ummqedsxXfJLqcdf8YWGS5tMK7M0nSuW2BS0SzhmT7u8GjIYoBoY+QgVAcEU6VWkEb+C87Np2My+
Xgj5renjXKvfzTqWf2TxMqF8iZan93rxtwZanWogNzikgbyZA1ux8AJetpp8WhVuuQ0Nhwb5kFzx
YwMEWVMj25wkqUpSpc7Zg1JleRth47UgkIZMaIlQDYmLVSiA0MFIsrZEizGlLZFeATFotEjT2JGS
QnIUxO31c1l5nSSlUUNsA7KM4ry579jFQBA6EAj6L3J6efOGO+cAU2jYZ7oG2TakfVe+b2YVx2hL
V60H+siN9TFVL/vEINCXNBaLv20fyXumsc0rqyBkyzwjzgvVNDzwjCC/VJeKWVm91p6C0wIo9vOc
2jiLdmFXEQETLf5FlHlAlVlQPYaHJbrDTw+GCLh4TTm3FJtmv2PrCImioidPeuG6bW+2xrPJqVFk
xS77Ts5G+6U5gGbCpqSP8ippGJPmt72rgUC1PDQBMgAIKWYZo1MD7uvh1vOWAxj/lHdHCWHBV3hR
zNst0KBjGbChwH5fBg0DWAtpMOD5a9B5YdQ9wj5DUV8a9Q2eVH8FYSMiX8mHKmaK8hGL/B8Dxdzm
1UOO4MxdIc6NpsOSN7sicVseKQ/FnFRZrkucn9gBnqnBGEvERIGlyM0XlhmwTpi6/IGgRUvMDLHD
/tp0p2hny9PKR9f1H+LLyVHQO6FctfJOPu+eM+xctevDx0YLJPfnUvAdbYWaan1uEzvbJEW/irE/
nsKlF+hqSzxviFeie7G5uS2ItxWoIET7Nu9G1zUc5pdPchtsscQ92Rjn3XzW6xzcIE5y5O195kGV
ECldY/b/0m3EG3piNRgDXB4TNYzfAKhIZoJ7HftkQja0GjQh3yr9TRC1+l2lQ54gMXImBAX8IZJQ
W7EA9CAHFOMFx/Ae53EGKqnS0WP1qI56SLMDV2wGvbjPZic//JXotEUl8QdycPsybukKXdEKqTnk
uquNlZGyG3jEYJoHoLM1Trw0OonNwl9byeRPl1XJ/LrjECU7+i4xZ4ZhAwtdJntAud/139QyISZb
ZvHpqmbnRMzm9KkAreGRlBHaLdQctZkrjm5UgXcp8eY/518RINlDTrN2VIe9ZwQVBLU76hdTU8mi
ZDyHOYPVqqD/Xjsd8bT4uwJ5FS/Bx7KSYO0m6ULlvhYYLSrMfzyBJQMC+sNQHoUFwdLxqTLHqI7h
E/vfF9gTmBPsts8LM99k+aU5xKbT+wpJHCz8IdZyPoYeqQ6iGel/bNRP/a4W5LW+Hn8mcdqmVEez
tOqDSjs0O0Y2j7EoOf73ZLspXcjQMu0e+E/suy8n6G8k+q3gze234iPncmcBq18avZVGxIuvvE00
hfExSut3EJBvINgw5c79Xd45dOgzHSOakrCyWtN9ODX1RrD+LAyDF7H2N+jmvbIwG/KSoxv5uWG+
ssLst2whgh8gW7h82Ocvpi/Kc8zP8qht9rF/UzbfDizc1UIDptkHMr8a3D0r8OyYndfNbBho9dal
C897oxHHNce8UrY8rCyNs0w7adN4DXcb7DVtm+BCeANDvPCrYvKLmUKJ2+8vsG610dN65q6VdXQj
oYp/jmY4/8pqCMBxLz1twUjOYfD5TKltXxn6/6Buq3xNyaNOjDbUNbFe4fe52+bzsyM7qkJF8nqK
JsqyOB/Xhv35/N/WON09xXvGbMgtpynq7vW3FH+Mujq+3Darmsgzm3wYUkcCZLydn8K1GGaMK8QX
FXiMrFB4MBxEmFKuOpbLemAxEZQD8NuPV9X/h0PupblqebsvUDN3ma9412ZTpK6WIVwYIZPgEeRk
HNyyhzqZuWfsBEoVIRTUw1ohwwDmth9twkS+QnyZf0asHqENIezY3vGvEllXd+NnksS+ihkbFhhM
td1ZTrCK810YYntSmlDuKU//DA7Og1V+IfMiM5qJQjS2a9Zcw2ybFHfE883PvPhD50asyTLGQAD3
iOIYuxCq6Z3pxy1nr4gRWeiI+0boQ9xGMVtg6ULFmjdv/CN9q5c/8Oaa/SRW0aTOGfQWwsje+bCa
UviW9QPkupIkeUimjy16hQmIWoQGX61L5lUcwdZ2ThzQdcrom1zL0V4gZfQzQ0z5rmjvra48SJ9i
DjEdkyWV++pAvc+6vpzSDKHKisgYDp240WucQVHWA0o95YfwSDf2cazHXrZ0+DjsIURUFKryxqcP
umy9xM2AdPbhWeaBAYqkqkROHTcD+OB6CfTPxbTN9Go6Fux2q2SWQFlIUH4LLe99sLr+QP1tkR08
L66EcWDOnCg62iYJn3ugoo7pSolLtwiMqUfQYTy6hrBkP16oa83ccW/PyMZHz/YKuE155jGFZXQq
9ZdVASfWxt0bX6vyDXIlZLAaMpgAKpObetcE2/83HSGNI5zwWz/IuWDDPtukjhm8YSV/+W5beDlp
atqB0Sul41EGfAm2FqvyZXyxFe1oBiGgxBweAJxMMEdeXMoJsONtryEkPSfG7uQbeegXG0u2qEXA
/Key8HzcJ76b6e/KzDvz5ZbD8BDbkhAXhwqFI8fydedeAVE+0MI6F/b6ifbPioZgA1+guznzXEPY
oOJ5IhxaNZn7h+v18X2BbX+hhZQ72AFxH4aTG5mZZTs0d3X8BXLJlIHhHnsG6rGyhDrmkcZSyv6a
CJWAXUpkNLiC++ftZU1Y1Wzn2gR4AFhnbq/OtrPHofroYTiuQs137QAT0Z/pzdJYM5KSombmfzWC
ZJU09emzGeAimrOBVyvuqdqIb6NFLadEripdhLTLNrlKxBWIrFpygZFIEUcdpcmVyqAK3NPv+kjU
mRm34UZESC/AEPxoYc0cMDFs5ngRrX3znXORX6kXj8lTvnGpBfXxB1OUg+Kl/T+JF5kS984iUOo6
YlMJB8QZvkwEqYCYoAMzYmrs9hYzB83aKwAIkgmehbT8bEro2qtHFJ9DA0C99MZobTkirxsWcxYz
8oJ/8JW81DKwbZ+wJYu5woXusl4EG2+LGJF46NYhtnSl2UJkwCneaxrJ040eHcVAxs7bFEN/5IUI
4aztX6GccI6dRTHIBdaMY782+Y6+K5MaLGhKHhsWPUFhzjf7MK8/tdgIk218HNTobJteIWywQEbE
RI9vRfsLHYtsRC+lsIWPHZjb02nNNxtR2RzzOLF/3OjBl1cvU21dBLq66IKFSxSv3HJy2ll/0Obf
yxMCinaaTnArlw4+DDZG+34GhzrXfdzddEF5whpHvy5DdddsIBgIssCQt2YvEZn5Vqy18wEJh5VK
KR6PZ01q3me3mArKEOqbJE5VXA2TirsIwcsvpHg1add0N0pZC3/580HR4oBh5mGyJuhPrYxR+7AM
/fgO8B2JsTJjDkCV7X/I+F5r1LOuuVGQIh4e2Hu5Tgmi1og+7qMmsAbxfxFl3Ggktgt5B43rfH6m
LhsZw7+9q+bgY48IfLoB4Y66XlyLcSNMuPgAKb3WJ40RsCMYsg/VlAWYjwCKAz28we+O/yTeg9hH
mtTsCyeIlkoHvOAco952+bI1kKGgoS3Cl2ezMPpzwENfaQ3rs8AdpwveIhVDdNk+wWsa1gnlyeOc
AiNti8fUPYBAvLjV+PZTB12BnGvWhrE3omrwvWHMd25lAAPd6w2DKItxcb1DbTSjpE4qlVLSHuo4
2UidytIy+9Ae1N6xJpr6B9tAeG3uS5cczf/xz9/3WvZJofNitzeLNa6jBr8sVmwrhYBR0bfBUhRO
CKk3SjvIOznxNGXhls7C+JJY26oGLncmiBFBvZn5LkiRJZ4wR27or5tt+f7F06QYlD6lro0OGmI+
LtFy/563lFmkgV/mV+LYInKf2q5OapEfgBvxs6N2rf7+dqVcDyz4MVJJ/vZfvUgLM+QqIkiLE4HT
Tl275rhaGgl4vvuJ8GSUJGSm9LT393prZNRwbuH/WNlwXS/Xqx1k0nIO0nsh+ny5QbDu71Swkx5+
TQK5uwRTtjaxXFhPF6cRGJSFqP5t+fkLC/UrQUM+RVSX1DxKnT3f+Ye/NLxiNtsoDtR+IKGfydd6
rMJQ4GGoQ43bG0zFVlq+2D4C6M0XdetWydDaJfCXmpXif3TAumnsEM5ltqpPTeUoJxHRrnq2E/vf
bTN2ZqahE7401OvcO6y+eKZLee0HARp875pxqlxgRYWs/oW5p6qINd59BH0M/mPw44IfCgGCZWf7
qpBarjNITbRq2d0wOnng3eZuyxyHkzlZ2uE0lCfQMWkm6ELiBYPX/nbPaT3168bDeJDMsrw4VJN9
iIiwKsmRVWkDDaI60h/PDldLnknKmyj6j2vnV1SLPDIeQIV3ZL8pIFUFA9zpxFqLKtvox2QH3YJ+
6LgR9bcnj7sprsLBFSZwstMjEA6TMuoHEQsnss0WEK5dB9KV69+qbCW1Gem2pgOpG5KW4NMIQXvM
dd8iGEq0Jhk85P3qPWSGll8IZJgRHS0KCSPQybfJUTyOpZwQAn0qv+h4/tJTFRQsIBtpfPUqCJaO
JNubPFCKfdOuZpi8tMy++8OtVfrySf+oBDxCcgJWRuxw8ErP6n37e5U+4oflMnFpbBsE3/a5CrFW
Bg1FAjKBTfO6VN8aEfvZ16stlaME4txWkDyno3ndO0NyMhTuzWPZiI7Z3YrZOGqGdz7/enAIrTUv
wH6D1ylBByIh4dZQ0ByVLXxT8YgbGQxP4ERBfu5iBjH6lih2+bWK1ndo90Ild/GJOxwRYt2/65Ez
zbyz6dpfngfIzwr3hoYR8Mix0zr4PKEArNy1C/DK7b/qN57AQWa6G74YjOSOZ969zH8AUeAgELbq
PTzuHqtn8HhqFRUYgXeZmbrC59k60ShQOyUk4SPoQKyGqMwNC9Lt0KLVGzodLEEHKtXzYJtCE576
579Z5L/0SbElotYS+VX46FKxwpQ4LhDemTLxnnTRGAFCSnNhgrRmQjNv7xeW7J1OSzaZ97nMuEqc
CtDpCHXq6jlkNZSFyttDMJiHZFiAgJx4bvvGw/pUoLlbikiPexa9VjSw6g8/vFrg1nNAxzwWvebR
h85NRJWVK6S1PzWaUSXr6tgaygpoTSVRDUuepF8+/q1z6mVmWsVsnWU8Mt/oVH66dGDQ2bafvNpm
qtauIylNbCowoYPKaXh6FX5ivpMag2P2yixokGGsP5M+EovDB0+HMGRIqYuxQkR9ieuHS3blgik/
MWBRVYA2u0bA7i4E5fYBhrgR4JLNILPrEV5dBsW6rP8ZZTU0b9oNjxYk3Catgzq8bPd6xoQSp1Lb
71fzROPSTYY03N18SQ2Tx7/uwHA97Q7iYR9Ks+LZnSIZjVaR4VdHf0nWAgs48QvJbAFEOFNJlMd/
GFgM672UShLt34tvvplgbDuVGGL3ZZj9CdAy58u1CXHF0hSXc51koOLvsuO/2gHflq1+Y1lMaKA2
aUUEaYzsFdTT38V6XIyC4iycTeKhw2F/B7CqBmq1o0r1pdHyHgsY1j8v1KcZtRIrI1/FMseyeAXd
d2Hu+nLVEmhRCVt62ES12dZg1lAKZtUi7G3zeMQIN2VZzpNnij8+EF30NLSeG/vEkEpYBO5BM2xC
CV8eaAVEAXFf5cJlNKRxnaTxWYYHBKVizL0LAv5wsc4Y/uT//+b8K0ay4mckfzOIh8C2CqP/D8Jn
opdK8PbuxpNsYMeox7Fjm61kUF7szDsQ8uGqUbOUjzvzlVJMAuH+HuQ1snlwSPDSOG3EMEzIhKz0
sbtNY3Phn/a9CDTFbdvQDewm4X1sazF22SOhxzeQaXME/apY9Dmk8Ez2UOORuLy7Ag8zLFV3Lpwz
5AwEgqWyGllX2Uii7IAooIHQR0f+4MSizwZ0ARMMcKgX7e8+Ph3eteOO8XfI9TyCB/5+2kGejiJz
eLAU0qY7BTLSOgZfsJzJ6BJ65eppaZ7/gJsebxodikc0ZzXxy9N1Ld66uhsru1eIuPxmZcHDqI/B
y1YFFIWzQcLwE5jAj99gmnEkF2jx4374sM+ePvaBdq2lZbxGSSOd17mhNHKh0dzwiPSerbLaCwnG
nBPJf9cyJRE+HBPAIwMBdfnw3TTLbCRstJ0E0CN1QQoVNaGdOiEWnE4LXovtKUT1hc5LiLmg5JL9
pcTGfkPb16j0tKVIUgPQlrKGt4NVCiFZK69fQR4DUv6QgyJQ0hD4Lrzr7dI47aoVQdsthCwomYOk
3BKLB3uITjs0da5mk7tyGJvOdON2cdUxzOtJmhsdven2qxXtj2XBWBHqxEj1vwA3oMa8cdGZ0KTS
FZlVr3FFBWKZQqa0wDFRNQBkcJkIV1Ah65oZEawizurpClD4lRlbaxIftVKdkhBQpjWJFYaKmYsH
a8gkiZy/MqVzoaMarpdLbm/SMP7NaiwAleWK+ej4nsA5L0f9Nf2y1JZ0duxXNeuSQRKhJRKAWDY/
NoMY75p66uBunYYeKM8dqu7yxZ3k/mibjRsCyKSG2NeLAFNWZRb9VZ3PKN2ZTzYsFX2yF3W5eql8
jE/25lZooX7LbQVRVj+UW8ef0hDz18rw/scZVyvbsTz8FwPY7HaRriWZwGIcI590v/Plcwne1JFC
xgnn90TOpT98b7VXowb73q8jGkoumsoNgXhGhEL81qC4+IpaYl5rUNdTSGbft5HFZ5+KU4jd6f2O
pZxmiD/4fTAWmqyf2Hu56XWHNJbt5RKJ3tZdAquj6EWiE9Zg0Xjv4iM4gdrrMWATHm4x++axfZdi
4utJLY+BHaSwOLeluwzCcy8vWSSN45d9dmHHy5Y442vD7Z8YSp3VN9RIOchdPkIus2pmh857SCsw
fOfom63lDzPST3/tiNeUFs3ZDkOATZYqpxyNZAEXKV6ojrVvV1gdzhe6Xgy7QsVoHmcRY8V2G+/2
xfjxuaabmF9eg/69kKu1mttQ3BaEYiGOuNKpNmSEqhDCX+anzQjfS2nbiqAzdv+7FR8yUR/ydeXM
PDgp97RAOjPgBBqez1veP3bLtWANVqFS72kFdCFdjGv49v3EYVx8wOS99ZiJ4GQdbbyZ5zB4Y2ec
Iy6Kynt0e2Gtb2AmP/IDOAcYR6DpdeCyV8hdUqROWG6WYWgrPSTqdEX2kMSevglXxGseFX3egDko
xb/9eMRwSJ74zZdMghceuznqj61pMiPSer7cFyf+zRedAADaDbyTQhZt/r3sBKPmLdoKXZ5D3Yrn
AlJqRfdB+cxcqt2ws2DhzH8lY/721hGRGhNEm0ssWFXBTrrl9NHzjcZuP9ZmkqZqra7Q2ljd4Fg3
Vs9JK2FPhVfW+5c5tJrjalN/u+cMTL/fmXEJbtssxXGquKh8GIjnIhWccPFE/Weq5g0vKkIYAnrc
3HiTV9ZJQ1oO6QV2XOOjnFnJs532jYOTLtqJRKgQ8OaqlEiXgL33JnhvOMez/p7Wi86Rvd1ZiUpT
3FHfiPjKMpfCnqbSOjYWODJOARAz0AmdlIqX03XWzJpXXbKg5xAOdfNerub+bXrXsYs3GCbn2dI9
TYAYcCGX6vlKjPjr/F+PGFNAbFkGW+GH37f0zUFFP/sd85UnmUMyOUgJdEtdjQM1i1/xJRJLLCJq
CvuiQAq4IBBBPkX+wY5aMiEJYyH0UTdB+Q5m1ImE+7YJedBJBh0J/lawO1jDXxv1a8nBcZ5/067j
qBcnwdKZ7qCd2O4KH6Y1rf8dUb0CsNXtB4ugMd1FoNw0whuR3ZAgM4rlbrejsO/OviYm50YjIIeb
Me65l6AfVoSEltzh+g5jgUpqmsrzj3L6mTsTgJ0LMQMiV3mn5ghdJKfELSRK+PB4/v/1qyVk4Dun
Re5qyHzhrvAVX2AQZJ26yaASEr+H/eKKU7b0WozPTbv0nne92oHK9+i9MCvvxiT0NXlZBpfYCD1b
7BJY1+geNsQJxmmPHQzeZ5EXAt8UPqvYsfYi3kf+UjsReV0UxiRorBBPDXggjHR6UiIXohK2Ifzd
BE5x9OMGcCiWzSiddTm9v21FjIOx07fAYeXhZ+wfl3PjEVOBQUCP96mv5Kd67fYJaZzbohEXmvS5
08scsa7UZPCyQXMuM1jy4X/fkx7QiTg//FzFQuTPk9VtY/4mn8kk6JYAVzY9NEP7VdMeKgUW6EAh
hlfHZZK4V40QAS7OQvixQdMgdnOcrE7YQpGcnE5dsMhuOmGxNCQ5Ajq+u2NWGjNaLySYnaarVPqx
M15gxEzpEEQ2oQXPiPdB2e1AAUZdBig15xFx+7t2lveD58TGhHDJ+kPDYuFVEYSBrNThtHZmbFbK
5KPNZLE6Y5qMANvPfdb4c6nPAtIF6Z/Bbrivr12NZL9pfa2E57cXUtYxXml01+VF3dRN5LlZukts
0j2IWOyjnEiUA9RvicNL14Tk2tpcukE5ON73WB3q32nHJQj0QNCgJpYucA992GLXRPIrzZl8fzeH
q15uowuDkDdv26xk9MQ+D0naym2DDjfzA/ZP29sKq//eeeSN6dAN6NcdcwL5KFtugpkCk3OUg4JK
iGr37aXmHY/VI1KNgMKikfYf+3cojpVlpdRzm3l5z1mFvECmVVupLRc1grx9vPpnF00mW9Uf87yX
ObT2mw+JrgLYYasqgmy7JQZb2CnYwKjr05lB/MbBgtcXHYmM+j3sW+v4VMw+PjikpkD8PYAIiXNj
EEwKYgPl/IDBYgaDkgyeLi41ThXWGLP4/4Ec0xqh/YCAl0ChGbMzhtilV0Bwj/hb+b3QqdnmB/i8
SLrr7d/OLGyUJhTeZ3mdhCyciG3Ikf/POvshw4+qruXsYSJBQCADdutwXzA/LqdfBU6wamKoGoOL
VIvelXMu/D0fMNODvIfFQL1LBtvCrvGHz8HVr4UDLwpa3hUue0peQavvIOLoDiLYgSwld4OTN7Pk
PGNmd8R5LwmeIPvpeJ0PSISMgKamaMMmzFWRnZEagiTd4P33i+9gJUXQ/UQomR0ESgl1WIJ9fFEb
7muhs89NEFuHrQu3W4qNDC+oBYoSsZuJs4EKeS8sZiiuF42BH/GLamKOCp4ArBfx+HmMjq+FBtVG
ymDPCjI6iU/RaYN0J/pwHpfOCTUFY5hnVPvvmOmcVT2jt8u8/vR+XmcKAkbAykn5orWZgMZKorse
v/Lau5Z67XspwIODyRWzQpwohVFHqSv9NGbLuRwyp6HlxXjOJfxYpgBK19Dg76a+ytJiD0/ZHaAZ
o4z9NcWlKhgIJl7sMpaN+OYe3zW1AI7YGfxBILlfvZddULaSHd6+XhnQi2+4/KWprx1sRNE3Xf4O
kjpfvTDRqJE//l4YeJZoD8wohAAQ0QnQqnDSWLCaASR7LCkRL9tCiY6fE1ZjGUXDK27dLrwb8eX+
c9DAfK2KaUXVHz3ru5Dq1twHRe4rTv/2kg0pIG+SqA3IuKw8e/bHaPV6kPEJUS8o7O8L5F/eAMbz
8moxQ/JXGIe2OWJ3S8b5vNUBQF4rNrqTQYbIUQSXF8fG0MPPRx3Z6s6VzcuUf9sMBLbbYOnmOFYa
50FLgiHRAap7BspJ/Ec4jo896SqSAdtKeB0k/TJsaRvsdFvZkbDp+/iM4F+HJBetrgQyKD4rwttN
eseQS7RtjjjuK18kKGOFORIGODErxq0DvfNfo8Wq6nORSBxpALESavJuaJrbomjnL/PUsgYW61dw
mW+TI9EvHZfHalDKJ0BYDjQz4ZtOyTLtHGbEJWBwhTa2vhow/sy5aBiayyCr/u6TqDW0YiQsUqUS
GCYc9YMMGGDExR/Bm9G8bRVLtx+2mxgMpphjUNLcWA4mk1gFjTTZTHsMAHAyl+k77sisHViddWsW
o3ueru8F6MMOqjVtORJZ4ml2EQ7i5D5aJfXncXsSGkhxn9j/poD4I+48QBrB7LNk/iLdS6SxGJGT
m0e9gLxpDi46lpEIJ+MHDLP9aaOtHme52Tf6Vp3/4HNvYuVeYn+Akpmbn6AxgGMsMnbzrKSf0z4H
MhFNoiqMkmN1nZ1rnJ2iSJ0WV+tmiG3Ncftl/XC/KExCmp2iwH6uvDz5OTl9k1hT714V+nJchyRK
sidIuU8ppFva2q/Ocxb68QuCWhCDB/pcVXSqN/IfJBH3ZRJOAOnHGsEUkvrmajOQy/WdV7aQ+7Zn
fMcRFhI1yR4L8mq+ZF340sxSXLsnu3FCa9ZJa2U4/bbCor/+e96wZxCecjh45TNM6hr5mtVworW8
PXLB+U9IAtqBySKI0oM2SGqv0Hrd7ZJnA1ro5fhJZ31eo2gXcv2UlJUEucfGWRPjPBdYjIhy8Aoi
rrdgaFu/ztXDFH61DENnZjNZQ+vsTnqHVXS1N5jTxEEBNiFiXwllXY1UOOzdYyIOCKZ+DqafQ9va
VeO7iiDCEChSqLAppqRn6Bw2t13w2R3b+8a3rOeRN+v9k7hhYJW86nWyK2SAmMSI42NCHJP0pErK
eTXG/nlenWn36QuFiW43a5M994EoZAsfEr2dsPifZln0BIskRR37slApGS79HCyjxStoMIYcij0V
da+UStppS1SUNo1fsZTXiwOxqtsLd7bQj0o1gLmzG48vlazGAgIkjVjDlXHTdhIJ8bmbdD/ZCbLF
SQfz+qB3OvJEs/9H+fFuhyeRh0cDpnDxXrhPREienmpHLqjMsTp1bK39ARxTewucLld7lAbAtomg
b4cXWn6e321p62HX2HZ/MRsNc9lb6ZXpAwdUn3s0a+iLwr/csjTVWnDbMPX3+70Xd4xvU8NDYEEg
qIzWxyHA3eRQvtAMuyHIpb9TYf4nCMz4heJIWlGNzfbDI0ZFtqJuaU01dSy+uB80r8hwW93jysUy
Veudfhg53r7BG4i0fODJAihTtR6h6pU8MKMKiZAdMtPPHfWZUoxZHz7Sdbn26LMobN/WS0S+s1dd
Ii2Z46vSlZ6toakI8FlygK1ufe9DMLfGGOqHjxljEtc73QcOtkiry7+s86sB4Tg9yKubcT81k7Cx
AzWq3E0Oyx4SAjCTBaI11qOIXHymV1bsF7+scDVLhMAMSzx/NxOzo0jjNW53MPQUw+iwCKj6PPNv
1L0+1U0Id6sn62aWUdjv/Fpgb4p2gLuofhIErT1457BaYkn7UkTXnIiJ9BHIi3sUKeHyxWyDi4lu
4PyL+jCLDKWAvhQLueCujuB1cL/KCbOtYeFtX9fTrxmIJKLGD1cYjVdSHENP01L+TqVCYLqJ1NBV
zizuCvQ51SRkw253gXwKdaWnT9a7ac0QLJ/VgvW9w7JZlMSSNinWU20UfLO9aHdrad4ocSPKEEr2
RS5d2beJfsc+63urLYGxdvBCtUM2rT/3exbezuqrcQ8M0VPELHBzgccFTCbmHJOZonLSQL+MKeD7
W2DniKNRJeBfuokLmWmTaYULsZywUYLctqgz3pkN/XgEoTA8+uPc0CCRuTrPaqBAkzTQm+Gwfb0/
YT7x8boCo0kpWcfWtQ/JWHUgOIwbhN9wODLIudFgn5Woq0aLWL0bvSK+dBnKEKvm6IqegtI9E8Va
bsJOghIHfD/c2vI7k1tPy7yuvIh24ba00Sae9oUSjOkkbAU4yzK48lvaiRqd+q2ABvW8pI6oXa5C
dmfVrQfTt0IhqbiwP0n5JRl3Db7/UUxfJaW/iHgFscTBDoWUU7QJ5ZOv6r38I6cZJJGbx3h4bL8s
1cCrKvvc3Suu+e1r4R3PkJg5j+lVzeHfQJtQv5bNfl8zKIjefK0ADSPtvFYPq/xyU6jlfSgduc+1
cN8a8u7j4BmlQUAPsqcvFuKFFi74ZGKTroOO2XRUg2Y1zh5X+HlofoTvTH2CjkrhgF4SbF7W/VqZ
WZTsoKm5P9fBijkMRxx/IiI1969vRgp7lYW3TYGOaSkIr2+u8F30Hwui6W8RAJv0EL7uav81p+KZ
/cx9GZi3FB1SQF5JvelsLXC+nuzUnAk9FvRst+iOvDjdne8LsBtO/M23H/hg9SbtpLHXDO5abe+Q
zQEt2v2CFnNvcrpf2V+0wxI7IyVytCSp6y7RtBB4G3I6iI12Rk+QnXeuon+WUQadywzB3U3m1MF/
TBA5UCRfZq/vL3KUKaETV3qD5G+Ey2+Q3b0LSMj63aRtsr0q5IYMSu/5+Y3d21/LhjEa2LYFY+3Y
wCnq3uN/XzkmFnx8kE3fEe2KIFL5WWid+7AmPC7yaKOmZD1I6tlXlnQ304CJUjKdkFPooGBz/Vdu
RDYdTTXATLcyfKcvJ/PDSB5Rv2znixsPBrpKlgs5Fsk1qYsrgUlcx34+9YKKohxsRSA4K4vjHgFc
HBfHodEjyDSzIe4dUy1JFiplFDvTXUfH29/l7J31z7SuRH56w10+evYCUGSbCsg/rrAqvZrsUH4X
rCHBX3xBk9E2lsg13ifwErTPGDh0JI3IEpJ4VVemEjmHimv0iKAP0W8soRv9pRg2vaj4abOzNDw2
MMXsaUOjrnt9429qGGqXolSwSGMTw3Ll6Zx4/LGfOXJ2jxz4MAvaU804cXFNIhhC5xA4lFXx/B1A
tVw7hROoqtUOUVoZ/1dkV1nXxsWVJ5dzwyhFbGLtFoPpzNLUQe/kKxGy8AHvtj4X/zJRPW+BBB7/
LKEWYDfAwApWXHdEfVnR2wZFoi1LMreYBIrUJw8odoxfrQdiWowWoPxkKI5te7MCvCGh7xxB6OT6
Wyb82RtSIBu0jW68Va2qSRclX09Fm3KCt/LZGtdDVouF3BCeezAL9qQEWReUMqN90Y8QBZK961Cw
S3MwXSBLqmaGft6pdWRJkcRin/S7448LmhkN9hCCLbPBR58LjQlcrogP2aMLbqGomfR4mOS/8euY
7AsreKuvQNW9PG3cewo/mhgSvLtOQTMLs8RbjCCWoMXRHsANAnUoC1eOBVOo4jPtljw/mwHRfjxt
LlukgdQVMmhpc4BP0zGABXcs0JDd/JlSUIHpbeH9bMYkum/mFpzF6/z7iklPw0c7hllRfrht+ipp
ITmWZbUvCV5agA0cqYwgHzaQZbDLRMbuPSjmVLwA3Y1G5b8P3nZHgj+I64u05NA+8NrbYhoD5rMX
39Fve3ZsG9R0Q8u50BWe+6Zi5XB5bDGfRIYgeK60ywBy83TIGR52XY3pJtukRFXUf1aIUn0O1oi0
nRbD3BuQWHsT+qF0wGi+HfWM3D/K0ZaYSN7pLaUOxpB4JNdj3xn8OUTlSliD2o3Zgy8CTJ3PFaMV
sZDc3fzZScAof5NTOcK499pnXre21MUB7rbj9It/Ih/J1XQK0Zs1Ltrbk8o9kFokBtwsZQG5jlBO
J+jRQXxZ576CU5xiUgjp6F1ys93PekyX+sjwdY7LNC5g64UcEFs/nFZWYM5y2wFEUKWIf67OjIoc
cYDAFVAZc4QQeQ210iyOrjoNbMFUT4BzM2ZS1m8g760s1bI0tx3yLo7Ue6bP1J9aftBChbl7eNwh
jiH0zUKXr9sBFiHB/vUmE8qh0rdhta9W53v+6FKCLWCUOKZI/BjCyHYWOvcsStYdkLJYHcqmBIoo
RkpMfCHBNr2Fy56n+ruyD5aIFseB4gGN3zw8/BMfPpSvOaemhU7tJJXyEPPCZUYaacr02uTOQS7Y
O3Lb/jbnMo0mIDmavaITJ69cZCCa9DhKTqzy8FrPODDaNU8VdbXt4LZ6x1IayKoEbUYH6Zh/ia/5
wUgQJyhnQ1T63MlLMeb9eouIdAZv/jYFlt76/SUDdT6Wf0sFNvY6nifXMDfcHMrrvJU4WXC9CH3C
eKZUNq+LLU/42FeJRtJc54JDbhigszmi7Cq7KRMlDZZwZeVuAvJF8XglL5EiCJfOVNZw2fYOhCgj
QJCZO/Y19MrCX7KNOZJt5I0CAalNbF0gh8amEjcSg0QSwwM7xIvCKHYM7cD7GKfFwmC+Pgf0/4SG
O/vFESn4gbiw8kj6zUa0BERy1S8jUNnBJIszRRvzuN4ecErJ38rpNFZL5B1noUxaG3kpSNWuXGxj
ejiLMQ4dGaY4z/QKQJSjq/kP9fiA2jWwCnYa2v4cYo+V812mLDOn08rGWX/E2axSHfeixeNsqAWt
OD3T3RPw5qykq4iB55Rzep7BxJcebhjSvPfQlp62bbZ9km94XjRfa+sBJD91QUoXS2tzaD2FxT0C
YCnulB1bfZ4aZ67XA+tsokVEP2MVuiJEuE1DPjjsAN3WdxZWCOuwhz6vbEi+ZZq83mN5AicN0ZSp
PXM2IOsxO/VS0MSYyq5UeMqTqY7+/1OWuU976rDILqgxSCWrJzAQeKCCs4w+d37fvKugnu8P0oQm
eEo2AmoORBU0AgitwLzdL7gD02grFPm5oWEND7gAmkfmN6iWLfgZX/Q2ceU4UqXvBMnG6j2Bmur5
ADKeO+yxbuhGNXQ02OyTbinsfc/sOQWftNQnNy/ZRC8lophXElqCtxV7/zorRYMQ0uhPXFhRt61w
qybpgE+pn/b7Tk/FzUq3+EY+QFdrPy7kQpUHxv5WwnlIEDaX5iudHmkCtMlPTXInBbuE1uaROJRg
IMvV7UdDqrL7NJUFKqv78S+Kx8gwpe2pd3Ho9BijmbO+ak03kvHFdCDdQyc0ObgeRKQv/91Fvgrb
ac27hKYyMRcC/gdhtM1sVArp4HREIPdWkKxBnDTUm49Yctrz7fwlh6Adnk1cfMa2VRjUIIZ3DwHi
+Re4KzfGzqu9hZI+yT2Ex61Ryh42Tx1FO2IRq6AeaMJi8Zpl52aQlxmd5FbyKnvwFwr7LH2KPW1V
w+sGCbd+xDBeuLwsTcW89SNtYtECoADAe+WuNTkFjgL1V8AsWdvq519e+8mSUzO3Eh5U2HjL13AY
Nnk4fiQy91Q0dLqZkIPKCtiJNU+tz1aQadtnj6lC45cWRGBq//OccnVptP2kyFpqt5myR9crxk6n
ZPvwpmZVIaa+t1MO1uy4KRDYKHRM+X4gM+iiQM2/u/8kuwR7EeAkoUJ9Gntf/IKpris3Pap/PljD
U/eiKGP6UyrH3xSU2cRGaf24tKRv7XdAO9azlClU38IAiiUGD4przJnVndPXSQ6uAkAzCm+Pi8jm
W+YRB1AhPzhkI3S2JJju+CayCvZVqYmupTQUKMPc6rahfNGN61Xv2y6xqLVDlTyJD4I5w4HuZPOx
5lKGWI55jxBnQ1CN4VnZdb5tyJUy5ijXwtBzX0L1BwBPasXoFaakD40+ZVBXiXJd5pgaxuEye342
JrVuLYJhPMfyc4yqAndF6dYcxEC8sy88qoxc/NxCWVh4x68OBs9yGI3XjvZ3s7ZcXUw4q5C3E80m
JPulVUwi+uxH4dUMCJBe/4sAnyVtOrwRgSZ7jy+dW8OD2+4G78yo4bIuHtbkOE2W6xkjDEEPMvKZ
5+TVHbrihAEfQT0wrYC0N0rBP0pcbDg70HPR0rb9ekJXQKRckTzDxtvbZmxY6pDcxL9JZG7V0Afy
A1yUenYlg/N3baI0cD8DMk3qtiP8pGVzA5QFmQ9X+WJT941DNwTXLHCV3KHy7rrVMq8kwAizLV03
upvlnottHzIydvchfynJphsV5gIXeo9tKMQ8h4R6fYJin4t9hkprgA7GNPbWTKcXb/QgNeuUOj8c
kXmu9sx1c7nt1SsD9neQs3SjKKEJxGgGLELL0eJ5Qp2eD6+jUHGADaFe0TiiH7InGeNc7FFKsmaA
YIm2vqj4adVcbsbi8FYDMxR5O6ni4pqUNrD//H4UKf8U0m26i5FXfI0UYQI872C/R+PgGK9laK13
kiQeSK0CKkaKntodk/MH6QeUyeO9+r74Iba3ORNQ28nfOVFHJbbca5JvcQE9dfQkqQT6HkO0uH9a
AFiNSbWyBdowtkCi1Us1ci9dv6hpeKYk7PnICEv+5MII1of6Oi7PY5Lk8rSSZga4x7PIxkImfjbA
9UdutHvF/4l/2FpA3IWUleFai9aJfpqLuUsFPDIIXLipQd35RcHqA7/ExORClKNH1tESNMfen/Zt
XxojNM4ucvgoPt0RA5BfdxHo/Lmm0rB1AFYgGfjRZgS0I2xtSr5A37CoMUYsJ37a1bBU70MmGt8P
NgG9XSPorj6NuvMzjCUDogFOdTxrp64Qk+06jSojuDvDVvvdwtN0RqeHvE88WpQk1rMgsNF2cDDH
SRNw/GiwS3tp4BVW5i0tMv8nveV9sxcrIQW7rYdan0DydEwZUBL6ax+JyTP8zPPWGFoXItHtJMew
O7tYdl60ABvkOvk9uF1gNU8WqdMN8F78pIwxXOOMyGIAbw7QN5TD33752htfhPx3n9Zo1vvRjpFn
r/cnEM+NIj0TdNDn8IFUJY8GjF5XUP76yIJ6GC6h9Oq5nJXwvfV6kF3Ts+Fszw4xQaHe1edb/t2H
2M4gkKPt/vcwMqnpJcb9LKKmckuZ9TeysmeWXJkxIXs6IJcWfYs8/iJRRNCHbF8KLSdq/vLK48od
CGPWaYEf61e3kjL7qs11n82J5ytiaSecXYXnsz1zcZOYe4SEUnHr+CdhKC2yLNEHiZ5mEEvhAw5m
kE8SwAAIR9BFtMVq9YPwUR/pnQu7IbFHJ60kkf6a7LTeDeTTOvAoDntMSxC6S7j6X64eoQxXW4TE
OwxPsiS0R8iLoz7VaumeJZK5DHgqn77zD1rrI8Wfkzu7HL9s0wBcVAAJ7yDn0TcRRjDm2XIvSEPp
ZW2aq3Vdkkmx3VfZPG0YVjsVlqdLguMbheDNVOd1mjoaRSFaehmft5Gm/D+fl1XvHhh44/fu1fgb
NfkJbYzajeMTBjSpbFwL0rkmwgWdVhOeW3aKkRkkUz3Y4i52DgRol8yNQSZhugmYFvKKzOhFBMYd
i0bxK7TYTWtxVL5E5A2jsClgyCjtJ/t7MUJxQ0NJ4TzI7XOwnswM3wnEQlHUUmluFyKbK8T1PCWD
Eq//Pl1yiUDV1wyDK1PLdO+v55LsB6PsNUVLm5rQkpE94n4I0/69C+U21nKkWP5XOkIUH9+ZTSDE
EegADmaIHWA/3m2/Qe6ZzLIHIR9JIMeoNw0xMjJ4wUP0L/HmMYJtv0a8qAu8TJBU0qheIfgSeg8J
6VDmNIhwNl1oUyBtcKs3+3He37HzoU6kwl3bgbyoECa8zeIVd+raeclFyuLyq2jsLByNI8Uf87Wy
f0zQPJEeP+qTVIp5d8c7FQ+yF7QFDCl6PR+r3XMFRnFAkZ2feAbVzGgbzBiPG4XS9oAfqNl6gBnF
/ZBjmEY6ofRS6OGVoeGciLmllwmVXyEVXn9VN7FNkOMxaO0zAnc/hVWpMVyUMo6g/Q5bOG8sP70k
zandWrRZxV9KzfHQPfIaCuOu+zPibO/aT6pGyVT6xCH8sz4YEDCdcvB9V/J/yqe9fXDqId+6rexl
z9zFcqNfLTm7EItcqvMzvwBnHqO+MKImDtjqVO5v7YWXyMfCTkUbrQXC8fu+qJu11k5y30G4RLkj
Ud3pRh0fO3GnCr3B9bpKFANqsyTMm3m4y3w/X6GHuUf1IR7wgWijpuktOnPAEizxpPeSz7E9y7WP
1VWhiZvpbzJxEPRSZRj/66ah3wOvjc2PYVxRvtxLKLrRG5a2nHFdVyHKHU/Mkkt/i874o8mwSNYP
fXBDT8iuV1QL5g1jW8EidOm7e7C+Crf/doCg3yXp93si2CO4Aesg66thFA56ALEpljGnuL+W3sj5
egHIEPacX+G3qFd6cLouUyUO1VUMzatJqlVjMxiVShRhWOyeJ6zRNYJQfSafiN5DJeesy2CWBS4p
TZcSaZ1pKEXfbmOyOU5kWiqazTBvH6nHkkjqBOl6CY/bffB12z8SjNH1aIdi4vM6ExWh/Sk61BBe
TES3TUI+M6PuR3jAEIwz0V4i2n5ubzBJxmQ8gl5OS1f+8PYAS5ipagX5AUqePGAuRrHGbdLG4eCZ
JafUZOxe+Zw8nURX/VITcfkzpxo2d/awO0xMy50oLQRzYC0RkAV5X+G1a1mswmf1agwS15rxVs14
TiVu9e40MqqOkDV5xDeojWD4twqt8NCaQ1JlZI9wOYLKKuo8E4Fsywh5yjJeUhjgmWd1dhnZktUb
4A0EyNgQq5FSavZUDWtGENNDzM5u14r6gcrRPdk3j5q5uWuSRlVwdEk069QrT2pwaJyxEqVcRd4y
9t4+eBqUlm9KmLE2OQqvmTesLDxF0k1PKXE1CSuJAszWsgQ03iDRrkQR9LpwENnr+4PfLAE+OGS0
JYBp0wyGUzFn4kO1wuyrBAHnpmBUWfahND4aranOcex6x2gjrjKSZDcAJqoK40cVIkSLM9RFSf16
Ytey++t4llO1yk4sitSSf5deEs61yNpurHrInoe5ceASVynBqJcfKF0ZtT8PPfs3IllNNdRpzHv3
aq0N8Ljeqc9auFmyPRda80ba523Yx96UG+PiubdXlGFr4U1D8Ta1CVyRYNuRTKLqK6eJcgH2UsNW
41pOeugtyp5ilnN8XwwuNy6iGOAZbvzi8C2WZQaPwq1VUsxKF3sowmNjZUqMXpzk/M/fk4dvT/eg
3nwg7Blz/83KLPkyJvXBrVzej9lySBq3QmCBa105Xu9Rf1jibGpCbsOdFv7zS78Qns1ieDCBNYp3
vJccMCCfU+LD1dwfnz2AtaEejl7ou32lFvxy0VWt/FSyvnF0uA7SopK1iMJf7RmfwMjUKsC7DGG+
/hthHYSBpvkykKpqwEeZ6Kb2iY6rIB0wdT5RaZIxuQ+EA8D4BTJdJeMcClf7eguAuWmA0H2d/u05
jycm9EEr4zU3umTjY5IgTRzKTFo5dKgBmlLCNKDu5WBxtp1vehH87HXMYe2TDJqNUsMzegJrxVTb
9xkHB9Jd1u2CiZEuJRtOkhPgwUUS9OKz7hFQDGF3b7/69arPPr6C9xSuAxx1gTMIkHko0yf4G32d
F4Qjf90ZDExIbankqwnumFdT42qtlLJV3Q0LBusIEpFEpCGMMmxxOMMzTHRWRPe+jQJpJrav1q2O
gGVKRtjDHd4n8Xkv/eYwX2PngNVtSvsjgOgncWmiIHMmLqUcwfR1hp5rlWRy5/zAMkZQYiMnc0PI
7Oir0MZxMDcLjOmEVWsHxKrL/4BVdtdyg7Wiyd+YlJN8WiP1f42q8mvpJUM0XxDRbeooPHy1tEV6
BrR42BYVP71OShaIg1DWspp19iV/28dEMtz4jb8Rj2lv7fpGTWmNPC6VBSCqjTlEDpCd92EsKem3
NHGEocR9WllBIF/ITPoGntvmGdpy+MyoJt3ee6lXt88VqZRbFVBTwvGJNHh3gclEeMFm0+7QeCiq
eZ/Px0Z9WcBYUOIkRYBZUcwkQ7Do++/bLomV/ToKKtPzQiAN0MxSCE67T2RTJa4/8YzuKjZYPJHS
/Ue8sBX57sk1nYbDMvYy9J4USh2m2I8UeWOeuz2Me6x1WjEO7lL3qFVucfIjD7R/C35Axa2oixIU
e6yrjobwc5sJ8w7IWqmNi/iDsb3zugQBMp518gKU5yMKrQwOyUKurmpzwbQX8q5HflWe9rpIGdaQ
vWnVy3jlBaubi4thEHuCIvy7QPvkON7qUf4kveeXdI7M7dFOdE2z0hs6es2nRWisNvE2/8+6zge7
old+UbE0uVM7JC7mfnCrhPHwJ9Z9xwU3sK3SDbnAwXleGNYMb5QJjeGB/MoqAR7oGmtQgrAT97rP
lkObM6mjuqPUjtR8HjmJS3mnv+Osv3hndGr3z5lXKQxN3VVdgNbIFHqDqZ4sh4Xmm16ZFaeUCZu2
knDLe80229vDQjA/Ve1Cr6Q9+1S/I8HTFOho8N56qC3OxMiEwyIq0artihpX9M6RzlHaksvUvc9o
+FVUQKJl8mC0mxST3RCxjOisPwZVFTOgFajv98/mxL7kav3c5dTFA47EXYiZkYg68f4zfdRw7RT+
ab+7OoomlgaKb19rHkKELTQVoy/x5/IOdZUJqO/XRwXgiP5BcFXRpUcPSC02ASsxL/eakqselZmn
P7CpjtXE1WTGFNWqTVXCR73Kh/uPfsl5c6BJj1uRFf2Epa+1EEj4HIk9gfE/oa6lwtWdGAiIn+NI
+H84bt2zgvDpbT//0/oTfBwLIY39MHPbsRvD7fTypS+Ywleyq1pvpqa1MCvV8sAagoxnXXOv8hAz
Ksl17kIcTVcqLY+adetq5mL1fkqLF7gpMBCSlTTaEEZ7uFp0yWBByZUPyvnBYwagGnbHFy9BncuK
MSmWuF9ZgRBYgc9CF7DxXn4os3swGlVwYA4o+WiR1Q5ZD9GnpXSAPkqQ5AQWBcixsZX5LVK1oHUT
ZbwWcNmlDC8QgHfYRpcS9I3OhDKD31yk9l0bDPFgBNCTItQAJcKztvYZq2hRUVQj7+1Ko6UnHy2d
fZchgz6ufb/NNuMywNumCnnST3LSp+wh3ytp849Fv97OV9jrT2yYzCZxuzP/W6lei0vskYaf7v0k
6FflUOAd2J6nJExlXSsCbTpkk1m2pW8BMZ4wu8R+pXTjJB9KmNKmbOu0GpksQnNUhvkKhUjXSmmC
pxdTIvm8QcZwL2uwVxfkUx9ep6Y4N6NfI8ATYXc2gj2Q/URsUXsvuTQJ0YdKkz2PyCEH8ovEfK3t
zZ2blBwj2GLYavIXRHSF5ZWQfYAlIKoLzP+Xwy+9X9DRi8soRye+VTSS7bt+7tmPpRmABv/SV1fQ
F9zVbDp1Pk5bwyUPxpJicTao9mh15rdzGkyB/Z64u9qN5JQXO1fQUapFIaat3nilv9+NHF4N7Jv+
wdqnjCcN0g0eSxnoP9+Dl2GH1KEB82/Z9mEqT1Pfzxdq68cYqJs5W4Z4eo+0UT+Nkw8zwyLWZ2z3
2sflORT2DUq/OgBOf0+AQIHXhtldytOA6l3Vw6LkvQnciknxBkO9J/iUzFFdQMeci8SUqWEX3zyM
OYBDJE1wMOn4x6ozLBEtGl1LSF1NRawnsrE5B6eCc/X9bwGrC+jCmDSiPpg3Q4EfB4yn/dB1Kgjc
DX/uKjLvl71dIsE8UFMuNuJSICQco6xbpWEjEkAm3JeQZPcfZn9eDk1iKO9HWRPDE8/eXfSIEJoy
OB7eD1CvMJtc1RZMndX2hyRmntOUVLnOX/2QXrLy4CF9xtzWBWEiLiQLQ0BiABiNNMus2fkbbUFr
BPOHoCyrw+FjL6r0bGgMXE4JOVM9zXKXs84s8HtWgnntsTZCRb2IsWL2oHathS/RuEI9u8xphpOe
vloQrKlwtmUpl9Ld2+AGXF0AfgD32OWqIbARrco+801xK3NYlGFhImee8q3oq0EB8AxFM5MujoGc
+6w0pzjziY3WG3jZFLxk6KHvu0MRCb949oyfT9K17KHYmgK7ZA+xtVokizrIqgHv6XHBgh9yKFaf
YYrtZobCDaLe5nwQS0gS0sjvA8mqtfGxBqfvEwadSPAGw3A2hZBYIBdMws6tzH0JOpfcs8imXXRY
D20cv5WbOjskGQPmytSyCMGj9eSgRtWsnzxgdx0OuuxIOAqS+dviu3diiA8bLMH+4k7EhTnOO4sd
sD4Hn79iWDD5ICg8EnoOqTngNBuFomoYsr23GUmBmtG8IF3AtpZd16KiolbzC38k9p7FtTymkPDR
aBHMTh7d0823nmZyrykWW0CG6FdRtfnIvaTWT05NMo5StqURj78cIgSngEg6eZXqnm6SD3bb23Ib
6N8lTsVWK4uUQ7DFRRRL/vqhG8Ko7MItWqkpfgZshQ+h6M5KvCTAPUqXAA9aKsdWY2+CKdvQgqAB
8yaZHDj5UaCmfgJcigeEYaTL6j/zA5MfbsMW9UoPO/RCgi4QBj12NMkX7aRw5i267JjD+blk4rlg
4wONurHRysOSsN9q4P/pmj/AU5DV7jwtgNIYnqGxZ7uohvvBBkH9cPMb3uFphskNB2GdHCFJd2Ks
wnsqCX6VPnzhzEhosJnmsmb/8jGFAsFAdZV7OAxgSYrMYD170jVepc1NUq7zyuLop+HiNYLIyKaf
kty2S8+vuOJIm4LjzNaBQaeqGoHD7oFGcRoQy59dsYQ2n/8phY8MXNutJZ70kba12taJSRPOVQpT
0NLNhTrarWf+OEXnomhtR3sFyS/W5b4BeRL6Pwh7yn78qew1FUR4NWOuTvjsPmlBSDzPnG0HW/Iz
hyAzY83BNQK8id/x7/DNKtD5pJ1FFCVj3szvHJ40+FtguhQ3hbIz6DNuGjc++egbIr+SMvjEvKZD
Uu2QZ2hzwRaK3nxUCPFbtobOsbpskSSHWWw0LEks/kMn22LTESl0YGrxsYqcqoBZHANy6xWWo/0J
sCD6Z26ZY6tc7nYS9fGpQoPpkT/uox2nuhsuj/M5wj1goSoJ0AfCaSdt9H7sV8yUzeRl9aLj9UMM
Kkw2A9ExsO9QqQBI7qQYv1oI8cD1OPwwU6ZqqcWJByposf4biexysY5YQ/SO7oSiIMVOXOAKxpP7
kyRBz/pgdwcWzsQPlaChGO+QUNU81ivz0K5vEqtiMpce3dZ/SagfSuZW7gDl2fD6bH7L/J4ZL+3j
xQ0NJ/Z7Fty16nNsZrYx4mSH/lyrcFRcpYGM1v0JCzrq2QTz+yy3qaJRqCZQ4okT972dpWc/XAOa
YOMYVuNtvQGLM/wPQ52dluvPh7HvrWRc+wwf5udwb7t0flwepD/mwxmVdOCaxqhZtoP5aush+Rob
l1WbRp5DgHIqxAm8EFm7lJgk8qtivFEAcb62ka5GI7dS1EHhVn5W1P1Qnt30hpmQTL2zXRn2zMvG
ruMTYjcutmEheaE4Ttyd6myyZxR9wourtMyddgEYtPrkU2VykXPZ8022oGmAQxHtXIx/Vi/DR5XH
CPTyaiQkx7FGhVgMo5Wid0/7tD5W1x2PCO5F4+t58Y8MhqfrzmfqNPgICyR87HNbS0crqD8EUUrQ
+aTIkscO+DcSm11OFtorxM6OphKnSExENzjWBkugy5+nBaH3vWngrgOzp0li/PMjEn72sBQ7NIit
UwtDsSrmftctxyQlHR2obXWnRMbHY/mERtHnxvZlG93KGDWmLyqrnAr9uQ5hXJSfZs7hrP6cHMRN
MeJuqvh649Lz5vzzsYDIbK4OxxYIm8R5akLWgHIhRsMLYFqNKphIY4KjzCRQ77vFyR0s2igosxcf
tfCVVWT7sYveo8N/DgXGZdeUetoLChbS2fKyDYOHZNpTAKH+P/dq0SCsEw2lY8N5/VNJRvS7NaHB
LeOkuRtUoE4MfeLkRfBqzG12FWFnx0V/et+H0xTvlMK4zz0YXkuWtVxlnmjoGksldih0+29CmEYO
7jg5RxOS7bnHPT4UkK53XoMdfV411MmdpfX0MMSZwYRqg9W1GY1GjRim6+MyQ/HdQ0EAqSYkX7fO
NWgqiMowF0YFezFllsRvt2KJfPfiIKBWpnwt1kJyIP4Vw36izIqfnhg87h8vx8MdNTdpnRipTNXx
30+05jWfSHuPrq3QckAFL/rLkSJDYPLzIeZjS4cmOytXc2vNNwPwakBa1BJ5/pyW/k+iig3sItlT
zXXxEeaE0v10ijwFj9sepgMFyE9gmhCu1dEysQus9oKpIGmM6vTAtRK9xJX6utF3jRZyar9dr4J/
a+EOw6NhI7YILzOroxR2xFajQm8SPE97YKXDr5BBjsO+X6ljdbss9uQ23yE5S7jh3I4NrVHC7o+o
0tUE7cP5PQSwo/t7esfbrmJE8I3zs9y/Ph5UiMFmq9NQ+f47i7ipW4bf1a5mQe+GOR6yC93SUoVA
sCbjc/wxuGU+yLPiB9xfeWc0uV7GBm6w6exV15/tsNuzRDgDbb0B6/QDhIRefEZpN8qz0wUpklWu
TYjlpSVQss+pULc7CGMRBhpnoBaDbfBrDtj5EoJpDRpF2iO0lz7BfULnD0x3+lWYAz0/sWhhEKU+
Hv354NSnzNNFoIXm5LJ5AaFyzDk4lUHJ+dySAOAJjj0N6N/9NTqg1yRYlyGwQqmx7vKaCo/Lt77c
3HnMel4zbIvcKShRvuJ6R+xYVqyq8ASvBzsGfEjNRb3XsyOYqF9u7VVTAGnaRB0ptGAR7pGIcrU8
5cW/sV9DMhNyezm0M4hEblaVpchNLEdtUWLpeEm6xPJ1bOhWJ8kQd7PdBhDvkal43cm6KuNgujkD
H+DRJOB5ATfWOfmT9Aa+hy2gXjm4W7zcRDW56d0mooZl2t8nq/krZ4Rvok06D9XARvWD4g2UyEiJ
4DujRvcEqfwB5dVJcFKgp78c7iuVfNSIeI6G/7ee28wCdOmUg1+hUk+6rOdiYb4VsQ6wG3jcpZe2
MhC9q2zZl4ndZ69fKin72KgQnLF2MVmf3yqQ6NygfSYMToCba6NOA5edr0zZ6+v4XOUus89UsbOb
yhX1Qk0msAH46Xap5xtUi/d8BwY0HPXPC+hSWuCQSuGcZR81i7Z+5DIuYm+FSUJygf871e7ICLAd
Mc7blHVQsJPBE0nG2e/3w3tgXECqR7JVeOz9K24YU/dNk3tnsZ3VZd2UyLZ0mL0Z6CEfvIEMGbNq
Qk4Iu55d5f70r6jFnCCNrOaO9rSRhHmFn86JmoBb4FVyZAVcHs2ofXhlqMUOEANI0mBWblioh10J
2/f7vIi8H1Aw5YidHsVKLzU72V1hhgVHHj/9F1c+kBOC14iwbznE+liTZKcQ/DnFeQGn374Svy+f
FFe0IT6q9oCptBWoJUfQeQiei/LPW/IE5xX0bd0EzvbaZtGA1sN/1iIrQ3D1ZZDvCQF0rOGLEj6X
bbk902tlMRveGaF0LrMWCAkOViP96g0BDALK/Bq54+yixr9B7kz52u6Csu3KZi6J7TJWM6R1etaz
OJo50VkrJFJ2c63Wl/jB0z2QwTbiMpGtuOiyMJua6zOA0Ni/HEKHCDUwmBCWDJywtl5TLldlzBGf
taTjGYMY+/AkBo4UvOjyyhl/u9NCPKdmT7mP0C8WaTb65FrZTK84xByaQkAZNZQjS7ouW8pGGkuR
mnhDFLeap/xU52EzyWJf+TefoDxhANyyiXFrfx/uaxFcGngs444gbUH6mAY+JHeTh5UTBabeqgNy
p9THFUwLnSoU11y//8yZpZErGjqXi7dvLI0oGgryRZ82h0wu3535N+vTTmXp4aLx7rtx6SmwP2rb
5TxSw2NkDhZMuwYXFR7wdzoDAJaFc9gfp+EV8Nb4pJaoby8aXCdMNgDkNRy3WfUJjvyUq/0R1SYU
4MljL/6y0HOJDBVj2EzXNhSkxYq5HOc2Xa/WvK3PtmoUrP2EcX4oBFvvVYtYZI55GY82Q3dcqUF2
+78ayrc6rmyQW1dVMcyflWq4AxRc9hk5yUQwSMQ+oNIABlh39qowbiy5eJ0b/VtxDcOhYdNkxUyy
ZFuv6PgfXPEmqcYLFrffM6g9evPbcbLy0AL3I5JA1SwKBf2KUVxEwtknGtDsAQAfgo3DKoGKkdZX
d0tkEy6aSvJdVk7yGl1OrN2Cr19IceMTn91QTLbn64LtWwAZs8iwGY0dPG0I/hxPz2nV0GDqYtVL
14mPsjFwbV/l2S98xTrMY1TbBugyRFaX3cSOcYCvbI341W+IFEktKgSoBBTvE2hVexg87Eeukbp+
uF0pObFZK+zZlswEXUr+BiK8B4JGGF6qCsaMvI2O2oNZRoFupemucyovU3MMOtrXzSqJo1hvfoQm
I2bX8VFxB2WmtPUpCqM5JSIBtpEIt4CeVIB2cBDwWkkYkRzG9Img/TPT4UBwts1LNr/9XosJuqAa
BfU2M4tQnjujEQT0uRgy1z4sr5jjfIlPBa3yCttwsT/1f+GE9WsAfUlIDxU/2myJyUAGE0ZNTmr9
sqhXo6kyN8+m8A79rdXYXrySaUDG9Lvy1o+ZuO6JcepbE5+dg4AdoySzBM8qs+JHRVRXKJ+kWHnV
pFt4/x9/bhsalTdRwdNnDaXNXOhuX3xWxCKjCSM0dSkmpYTEJcUzNkEVbG4UIFS/92qekBWe9IHB
eJXpv28TeCqY1NkKp/3C3SCbmO8RBVPHzzXxuYRqHqBJF/nCVm90INprv/9CJ9iT+xfpmqW7P5qn
0kwfSR/22e75P8uCnqsh0N/spVb0ShEP9bqQfTQh2apuyqiEAv9jYlwaemhHtutqI+3ZHHORjk5r
pN2+cKdu29G+EVBykDK0uTsAZ7/8jrAKs6bB7cbFgvVRid5EczA/1aVmDAmogMjouqCJ3bK+85io
260GdUeoVw3q8A7Blvp7CC9d+6u3TunzeUPZsVGHKqu73tPMD9kThTsxWqOOYQ/r8FZWSWCp3TSI
7X4SBD66IDqUqpWxJir9OXb2M3EJowB98A+EmWN2QoPcwJKlwW/Gt5PSfnGq6F3m4Ac+eRBuBwFS
Wr6b6mPRvqMAYUBmNiMIQDEksRoA2XCMJBEVdfXNK9oe+HG7M/6xzW8qGnQEUzCi5ECMjYIGuKEM
9NTX2LWAlaAJD+4wcpSDPux52Z978u4zU+kpSOj4QbdnHQTNybKW0lQboRT6OoRhlDEWxR/iMCI/
Pi6nGxCcYQkJs2qqtFEIgnf8Qq0fBHi+eh2x7yF2ABq4rXrYV4tLUbLe8BCxAnU8Km51oGnyCUIH
02HsfbYR1le4lLFR+bhui7qCm6Bcp5wVEZoZclWhEyD7DK/QJpQA95H3ljqILWIPaMsnCqaIOK6h
PtZ+7vQUr7qMnftdHwcXTKlHXJUWngoCATtYx1omQjqmx4y5gM9pzdLpBApy16Bjw2adBZ8scFBt
ugeRPCCIdVTRlZW6ntJZqOxujkq/pAy5QW86+vqFaDzv1XTXDswPAJ0Ld6Wz7WRC6H4T6Z8CL2rK
78tZkYoZksfj4dhvUB8njNBi42zgjPwCLq0Y1MDnObZU9W6Jt3IbaDToTRU4cmse6vGpSCXrSSKa
P/JcsQd4FecNHYQ7/mUkIwjBmtF7vh0/VKCJhMjhLiW6u6QEnQLAxkD7jZsrdNVwwHElRwKmBGd5
z6A8WJ/RMkSEeiSs7XHjJIJ5E469eRRw0QNvyxF5zIucW4z1NxHWdnntWOhDdDHL5S4PPiWMWiYu
EcJDCxXtD7j5l9yY40p9Hb1QcHonQTJH1/PEfBpK0f0gBukVpNUECH1wB2AwQB97ir5npAAdIuPt
AguaP/TyfSPrUcW/r3ZF62QBoMDb8g6rBSl3eZg5FXk03FJXe9rjL4omEYOsS1sCoD4vqCkQNnMF
P6fw8xAha5D5HDv92YKTP2MirH0mOGMVRhVtDK8enUErN4NEKacrs9+kt9kuM5aFnObmschxTtUo
qKrpNwmMRQIaxqV9sbHGsizDJMB40FPYucHGo6ZgLVSKlfueW9T50XgfjiWGxMgQOLBogPrZn0KB
nkbVway5c0XhvCrj37Q6kJQP6RghCSa1dbuCaXvcaiNQesXmaZs+IsgqNLOkl9d+pUpdh0ZG3Fks
ZhSyU4XPL4ix9mMyQIfkx9y6yh+kN51ViE5DEI7vDYaR7V4r+lFpdusYNpdZ72mUA44+4NZhREHM
3TyKKMpcCCQ/cPygCSjK4sK9/iLtz8kKy2gEEqyRQh71dl0tscxgUe89th6E2e09XuhccwqAbvzl
rsiSnC8rQy1Z5DNriT8Jy21k6OwKNtYlg6oPkJ7BL7SkjnAg8kXiS+7LSoMvVaQpBuqzpUwWSK2w
mwgQRDCJN84dRKrtl+VG7NYYM1QyRERYhg8GBzCV4IkclkrmdPUrQaLfu8Jha4uru3bEwifNUXX+
Zn6IWQoelgX98SDjD8UwyRxQJ7I8GoQwiunowhink0oG+AUazfutQ4eS58koXYMiYA873DlD6tLQ
pYv+v+EyVhx+5sDPA4mPN0xa4T1rKmWegFxdnDSAdjrvhqugpydHIrWn6exsdlbSZqZzzINr0CN3
QyaNFnsNJCH4S4Qx7ukr4aQ7PqothYmWV9GD7j+utRzMz3XaXjPYsjsOhH18n6HXCygx2lmVV14z
jCbrd1vBuwbjJjFZB4s0nJ3pPVxvOdGi2ATgbeJ8sb2v5u6NLrvtz0sIAnBwcKRlMb/v5id9m7O6
HsGipEtPjtwZu9GygyoyLR/qP8S+vFdKEFIn0zF1LMWtDKfEVrB0/yOlHs3SLDe06nLER6pHGRR4
OEdHWRBN/vD8M1opYr8ohVGIJNPF0futzcsvfUThzPXC89TmyD2tUIv2QXSiUmylScRt2A9WWpYu
GgR/DX217sdl/KstS0Ukv6S/87pyVABz5JmGXdXYa/0atQL00HWjPUcRwgT9DYZDkPQXlfTZ60F3
z8fjSMBrcp9iqPiCU5OxcQwbPryZoNCI6GEYhTNTWJBuua1I4mKLtOVc7tb3QGYtXq2IcgR54ceC
/3bOHwnIZpgtKi49LUwRWhw4tJfNsMgl2sELemkf4UJZFQr0olG4yLu0sBWoyTCovX6EFt/BWQAS
as3psvY31obYwzjJf2eUuJX8fMq3UmyUzfr2VwIXlShRaQpgfxMW5NMj8R5oJDLeHrlP23HJ0HiC
Ivr7tqX8x7o7A32st01nZYi31dlsr5YUZBP+74A8ft39xtCT+e4ZqBf2uZsqGJyTADN3gpvJYtDX
KpRxU5w9AdLUZBxDAciwFx/EaAebUun7sNkmRH+3CmNgfM7YU3bdamcC4ivFVgdtxhu0HzIVCSN2
8e0N88F/JBowJWdanroaiFGxWYxC+Ef6EPiFb5+RPJiS9PuYRKGlVGlqbV3CUxpugTqPLFPOWCdZ
at0OJJ6M7hM/4fX5Evo4vSGmC9VkYk32Wn2wEy/YUCU7+f8UYYUoTsnfjOWaU0GgDknZEyhFNO6Y
MWFLxIptppG/BOlWZ57CpeB9pT1FMBFC7QC7xrHmXhqPXwLDUhql84mDQ6kJV7A6IUnEwcNrqRkf
JMa8XDahX8Oa51uiAfIBA4JUw6S9MNpR0fXspixauOj2veAlDw3uVyOpd5HE3mX6YNBbH6YYIsLf
Ng0MEkdRtONwhvZwHvFNKCAUmE/brDmMgN+U9O13SXqm/plm4Z/Dv7eKy1ZRhqPgGgvOYIItAF0l
O4tXRp/b1OXU57+eeLPKk6gjcw11EhkgBdgOJj8yzWh+9lxZcouwxC4Skzimf73ACEq8ZKOPyHH6
uRWhgI4wjo24bE/voZSpfsXWGk85kxq58h1op+RYUR4jIh7OdfZjzFGD/ZhEtlpG1KmWp0wTDe53
KIp6ptowmUBw++se7ti15+FW4TCDOHn0L+d4DSiKt49CaqvMLQF4A1CPSQ/OQPXupda9cdleS7+4
nf+kynwwRS+A2/uUKvCMb/LX9Ms1Bm3DJYbO0xU73n4SyTYV3yTBUN46v8PhtxT8qz1z80xrSNyJ
qV97nHbOywxxGxeDPqssnAYZTyRgch9ztyzZXRxiwR7DHMGY5+a/DBOMFtJKS5s47W1z1jqp5Tnq
eeFVShVhJtcBcbgUYker6J+DDwHVTeLfKWW9jM3rH8OwaCz7aJv7PdoCNdx68zzUjZUW4dOIqZDK
dTrVH5oq75gjQRBJXAWU0pXXJL9p2vhcLLKY1L6VfNJSAcSibHEX1Gx1VbKxK3WGKYSD9e9XLNSB
NwQ8O00pot2pR5EE9RNdKCwRdMHsWsGroQx37KzJKqqBjo8E5247UBiRpirz1NO7olMBw9wMMpgh
DOKm0x+SjGQBEAo+ZteBWkG1o3X6/aJ3TzOPiStauaxrdF4FuQ91RPlf14NMbJ6hE3/hO1pWYATc
H27a9y4kGMFoOvf4kwPvIwe2DDQz8Jff2fXPdaKw1G9P9PKYPTtYdTKZqPVfQZiajYe77dp8rhdY
2MnrFmtHu5pTVlM+CHGBN1IH5nb8C3kx0CnQgfahFKPNq2qryRcZ2Q/p9vwJO3dJF9EfUPy0k03o
rdU2nECl8qHeO2z7AiCLWpZ4nDRciaR8FmtuRtYYH8Kv8xEF2/lRMTTbZLUqGUNiV6oirWM3IWq/
3j4bEnUTJxAlJIAxCoZptD9ROXkW2Ct2ZaFJ7B7v0zAWhK5Ap0qD48jfXajP6C7Tur2/nJX85ITl
iC4Q4pSKK/ffhhZ2rPq/hBgv1fcJQPc2ssMKidZBRyotm00HjxZnu/6skZ4eqzcr9Q4QnMEcKcDI
z+K8jvNdWbNSnFJDPOJ0R660AP4kRbTg/M1F7xG5pyYfvy0MBhBS0R9KUhWQhmFseueNiqMxRsbz
DtvJ4eZHzlf3uRkISZSihRRMEBL8p7zboVzmvXMnulihjYuavwiTIRkQDbDDruq7XRuYVFQfnHbB
5fNU4DtZZ6fOqpyWl/L2JdIJsPQiG/BCJZ+XpKDyFGHptXGzZNjVyt9DyDsM20eVlywmUOVGrIVS
aobCAt2NnplLjElB0VHLkxLdQ+3t7/fWBdhZn9L8erFhN6K5s7U4+6vdqvPbJKvlv8kif42RPwno
o5Bt3rYGwMcX1WoXHHXD9bF1EZ2/N9tK0heDGliP4oowyD6wW51VjFuZ5EvrlrGexo0BIlErvmAr
2v4T1+3tBAppcq0l+qWWceHPAMoPh9U5FUBmw6l7suaCZdaq/MqWD7tHdMNWYeeezRuOluou3Aly
d2B25DYuW69tGmPMRyhiD1ISDZP2ZhYGe6XrmgzOPywK/nXqFI/YKkSms/DVXUqALzTTwErHinIm
FrRtDn0koHoi0wNZAHx6JzCXgkoqd1j2ZW58lLwVx+z6ACt2bhFuMGvbZZcmQGz66+53zxKakQUb
avLPimPl7JlU0jpHCqaMJk1DV6oTU2rG5z0Phq6RdsTQjygpqkx22kyu6jW3ZAr/+G1l3SaqOPqu
GJn2FDnLIxezcbUXk76b2J4MFnopkbKR0SIGCkFEMsfAJ2yhGQ7buBDk9anr1WbAXMUXL+4YJBTh
XEWs44mNj12RL3pfkI+YGvzDyJfmI9QRabZ4+zGR5SVEVziafvZ0BToH+L7hSeSZ08mOBdQDUqRP
Fz9mF4TOgGzKnoiiFwQAKCThhv0Xoc20i+OaOi5b66bDtaDtFBp1lOM6sMFBsN7uufXab2VMAd7x
hUIRul3IFnFRChS7mENxgMNPmtu3B8f2tg6SXuTgpR5/BhR3i4EtXuQj4p59T1AwSy34AZQGBoTM
Ji6TGJ9Ob2dOP85WO5HG9eQGThQliftQDKFDF8N4IMZAepwaz88N/Yj7MOEC1CzYAmRnf1Gcb1wD
MFAT3z1MzSNr4WMbSLb9W+V/QrrK02K1Bb/zWeLv6dJA4AYWMWrMHTjpdpYto6k123tmbcag2LJq
iR5wfKaBT9F+c/Hg/ipwmzWrOnk8iKWbPRnd22hWp8upUaTOzZ0qtOVZ7CDhGZZ3oEdVO4LmjTcS
uaWUsNaTXgAQOY0blX/kRyksctfE28+FCs8NytCwqGU7hgcArCGYpxKn5/Au+0ou9hI6fzUXJMCA
EuOrQ1D+MyM7/wk1VL75PEEPoJaxBNmcFzHVgFPSLRDgrTHGQ/dqbp9YAJ5M4VRPEep1oa2IMtMX
I9PLowFgvL1c1gZn9jaHVPBbzab1KYl7mU9OaNf4FoSgDdJ960qoHgQvKKWq1lnzCKuMrgBk4kIG
Xo2vpgiFiDW7aU3RfwbRqGz81qvLwGbWZ3zF13FR37VZYzYg7YhKMzbFtB8TY0PUW1Nmkc8hYtGz
Ovgwq+ueR5Tos5FMGeSgK8QVGlvZdqUYuXMXhfHKcVGgR7ciPzaIcH8uXizVdn0K9n0F8Y/3OBoj
hozgjYMCW1M5u4z+3/xibOwE3uoFfBXeDKlmh77mbvnrepNV2iVHyd/s5PgwZWA5RsZtjd9SqQ1t
cZTrx7pKa2lsEUZDQMem7atcFvawbhUk8wFd8dBNpvaDj0ZCkuMkwO29S15RMo/hSnggi1iN4gow
S9kGjiUEl1QPJuKs2r5mvia1/2bo0lgpA+ZbBD2Zed5GOGCbsooljcGgB+d4uH2/yKOGHq5zn6eJ
70mIf1R+C9I2Z+RNq5DIJ6qWDcLVCBPvpCGvpwr/3bZMXuO8t8Ar/w5zMDe70wLZghmvHS3kPzYA
Wqad++2+9j5tGQI9FZzWioTtmO6Rdfhf5ySPfff583qxuIdAm3gmbFubeSXpg6pendvQWG6Ni3m4
RwNQht/TkFvFrZH+xBm2WOfreDyzkXX94IXb9CqXiiilpPG3GY5dJAVIe5qgwQ3OEHdtytqs9mdz
/rbycCiUXn94hDpTBWYa+snlazQ1pzxMQ4foyg4G0Dveo9bI4Sg1QVp9z0VJWgPOVDTyNspQIabM
rOPTjZJ4P4WkMnKkxO9LbBrNoNwabVLqo9m2yeinMMGMqN7nfLXeq6llN/VRAbhSTzmdmsH9QNHv
A68Og9R2RSuv6GhLxHQovJs1dcKNFslavUhvZf+B2Wr8lr3dY5h32pTjc4unkMEIGHnV3We81lE1
i25TyBm+2ad2N8Ugs2cWgCrsRVRoygEH5pWHBg2GT3joz7l4Swuu7X0dZcznBlUuUJKfWeD7Z2Wr
VyuOP6F8gfFjB2hTGkg1tyPbRF4Sc7iGSyHvlCpCaeYirEmX8f6jc93PXKBZL8JMSYJa40rvNf70
i1PS8SgvDoZioUZnAyGMy8FmExUw6oU/J1puRXpJ/aM7/fuikyVX2VwgLZcGgnryFtcHAufcKxoK
ng7cW9pWXtDtk9itSyAQJIL8rjhaUluBeNV9VjWi5fDo2k3kQb5aw1y1Sx9tRDvd2mvHLvXpVSle
pqjGpYz1j0ajcHhNyay9JlpQaD7BqhMeD1s6jAQIFrdy0NXa+3jkOJi8WWReIvNFmDFOUbwu308S
6m5B0EptE+yQoMqiNFOJfkiRVW59K7qwljYGawM9K+LbH1TJj4BBoKn9v1uvg2xCcLoWQP52mOy1
ppFv3Oem20B3VQqE9+pIh/RgxUGnsUK4scW8z7BXrR5esZ0SksVjEeOP3ED8J8+KJNjcyE6Lp9Vj
Pd7LFjKJMzKOyfBtlALySYxC33xnpwvTl+0GnYPRw8x4gGXFGRS72ShAQ2DD+jLyLDP7A/ovhJ1U
yfZggoxkOX3TfJUzc7yGkyKHZVPj4eX/Mzyopsr23jJjY9QWFeIgMlXBVgWfddL9kcp8PfI2dsiu
h/rHrlQCPcfSVRcvXR+vm/avUruu0uugbW5NNTHpinSq4OoaaoZ6K1PcMIEjewk9S4xU5Egr3TVQ
om0zxFCVIfpgjjzkhS+sk3kln8+qnOaI9OtrRjnjyECiWRD4n2wcdjxfP0h9A47joROu2hgsP7AF
QBDO4mGgAYF1P21mhG15Nre27cyOr2IvZGs6xLytzFNkbZ7y6cbTHO0n9lgQIXmcRjgr5f6JdNZ/
KYYh241/RYqO0fmHohu0CIZOdxBQhbKDVbZtpVQFhLJ5QVyhe2h+TDX46ocXkbo7cpfyQZdmlRW9
O44vXwlfKUiisQ0ntcJOhkiGLtBHh9BQt3iZ7l5sj5lgEKP3/r62i3sKN+aqovUHVF5Hdp8XBfDg
NDAEHonxO2UBAwbxdxd6rdLzN8X6vsz03rcG3bEINzrZHp9wEmjxd3g93SLfxTqLYqSbFCO54662
Xt9EIfy8+k8xMiJpAtJkTw2LnPlWzXoNXpaU1EwV958KSe4hBi2l+OUh90lGffjH3KuEh8cfY+mL
L0rswOBKU4/ByMXvCkdFALMrVCNzfg338C+G+1+MAyTSIWvgFw+HbQrHV/EACKGNEfTAP9Z6cJ88
yQITJE9CNqSSI8S90u7GZaF6eAtBnjGeXGBwzR/TajhecyKUZgM8nQojZ3TIsUlaua1q5goTNMQt
uj5nskOdJ2C2QviCqwKPZwf+3HBbr52WQzo002EUmQHm0TXrlomk0HF5hhK6g7hslI12BoCFw8Y5
87MBLNEl2StvRjoLrRrXWzzTawZL3d8WptSXlhhLmMrpsKpAPms6Wrhhs6+HtUL1IXbHbof8I5ao
5o1INzxkqi8vcXw8VGNiJ//EZ2z1owJvkWIs99nOsNKA/HDf8H62vhf+uufooaBD8T//Oj91aFqd
L1v6Mwagby4BamF+3dYkE11W+vcmsNeFzVpJlcMy9JXWW/LYCL+rbcAX3Igk0xQhKkGidBDYKKj1
O2qwmOfKmlQX9rsC9s2zflsezN8nVxfzHT2rr6yjFx9jD/H0HHE11XK2S+NZjMuX94Hoebo5yxZZ
IPV7eO2y6D5soY05Xk3Rk5BlPNWpkrvH1OlM9OPO2Nuulu1vzO8839qgs8ZyBzxm5+f8n3Qn2Gsa
/83dFXQoBxnQVkYzQeOjzYUIIbaKlQxoFVgZzjJ48CJ5shaAxVyCnZiPASs7We08g7EClW6xwb84
wQu33aahzrJ3FEtH47YFiQz7l9z++y8D2l7uhqIEFhDTAmmFfX2h/UQj5kjqMgYaSr7RldtlHHl/
dZHzOGOs1p8qUjTvO3FYO5vSmuS9h9fKRBWxAkQf3UfHx08VtVCgeRorythVPoPKjDlpvVNgWTKK
vhP3kVEwaAFVMeWRdVYHBefREHGwgxhulc+axWiLJP54rCuKlf79ZdCm+7QxF3MPqCHnzSm9a5CL
F8pxXGZ7d6YPQ+f4Fsk71xbJE/u7KbLxwTb5l8NEPCCLfkZGrUjDxFULZifsLVTCZhHlPuoh4Lzy
+hB+0VlEAQGTcYVt/FdjrFU+LgKPN4pcNuBzWBX4idXlkuR0XdUQAt9Tba7HIPwtFUHEiDJaBtg7
MFfq4V1EvkMu9h3sCX6llihIrVQ4JXx2+6UF94nTzbHUQAzCqh93eD2iEuJohJVTCbGXlM96Pua/
94S1WY2otNUsq4DuJFJKqpr0lPm0G96bUcDAZzj9qzEd2l5LdVFOwFyqNZnVyv23WiKkBD/IowVk
DB4uU7RbQtyXwtu6zB5wBWp2OReXg1lwa9xrNP6kUF943dYVVBLhNocP2FrZO+3FJt2qwPxftyaa
uOtB4SQabJ2C+Zen5wYN2eF1w/wxxie9Poxi+rRlhH0k0DKTTocFnKykPGgR66iYzdANdaYZtNqf
exK/b4FKer06FSaSDIhLwc3z2o2fXsCEexnQ0nIB3gxtxC2VZpfaidn93Jyb7UDgGT3cqreMEAAt
x8rczQzuoOk8SdMd7xvaZRNQJ0HoKrqoNrRX5YGBpkepzhJ9WFcDxvOgoRukFImwyIQ1rVqezGAs
UeAYDyxIELQWz4kt3HRTxLxrFcHPMpT8UIat8PhDdBBZpoVyhnDpCBlngPXItLQ0fCBjUzAU50VR
8Mo2M2h8kQ/+wjfOOctByyiglZchqJBNX8wb5e2wdz0R0yjLREs7xA+x2krVif98YUE68dpdwe+f
9i6c8fW4dvMXE07smuJACyBrJOEEYhhERwbTCzRTzqlCI35eRAZLFjBpdcpt8nMR+lroAEKIkfoF
SSwK4xrPIM/7YktJ+SV5OKNKIUUYmAcvHAY1jGQK00smeD3ElF3WuDSkow/wrQ8HpGTX9zmUlJOn
66JS9Ki5egxHDf1J2XyCvqH75CKWhIBtFIR6BYUcmgibXsY1H+CSvDGUb4TayKX+fIeW2LWjUs5N
Y1rj0298kxL8Ato/qI1siM9m4jiuhyoc8qnl43kfrPFiWo7a9XVazU0gme7bvUPiJ6ltLyD+VXMu
0cMLyEhJJxC4o9/UjZknpiy8vibQKJbHi0tVeFeX0XX78h4Zsi5U3GmwqHsp+aWS+Quj0yNGSa1A
FmVmWVXLKyoqoiB5xW2aoDGDcRjt/h6flTkLEKsITiQ9BF4L5bXsA5p9hnxyxWQP/e+pbM5TcBPl
R/ZD9xBtH+ThtPUzeLK/Es1O7EWpzV8bOIYIaQgGMr8Owjm/0nuVUGcdRdUxynbFA8zw3bqpkFIf
f9qJSIOAjh1i8cxXiyAeLBkMSpROwAdTqeOiRKJ2JNzLojBw322c1MK+WSO0fGRUytNre5vRZbmm
+ZajURXVSf6+rbH0kyUOXTwf2wPu66A23CP3xGX50EKwksdAWUA0onCJbYzGNc90WZT8D1SQPXKO
0eEI4PkPeKHpuNRTIyEKWUTo04BTFNOikRNOd3mRaV95PV3PULF51/ifUecnlxUzw71fGFS64kkc
aW/VU2L7ba+jvrwVhQl+9qybceXhsGk9mlfB+KKSMJSchM6xlMGTJeSp9PZOcj5P7qXyxTB7gbqH
oJGIrgUh2tKlgPJXXU95kYlTmMnuwjQeWiHp+UEfe+foDDgfdtH5zqBbXcobpz2D8d8eKqlSdRsI
whFpXYB/Cn9wYDCzJNO27lzCqPJ1BwOf0Q+BPRz/K6ZR4Ub23QuTW1wUxaLNleqGNLge5WSHu8qe
pKKe8qGA1Lxv3CAHBQGDq07Oh7xjoWd5y+nnK51fXcgPmyY0ib69/vdyBmaIAfMVf/3umDJy1Lc1
QDBScuKbuYpPmoIfZli1vNhcPFdR9+lW/ua1Tij0XXm4WQrkFzW2D9CxZURX+wFUU6D9Yx9zh6+i
Q+xDsrA/YzSmTIDWPxxqA6+3IFuV5al1nTEyniv324Nmp/4+tSW6UyCAUBuN+AmvdKIEF7kGa4cr
Dxf34MJuGucs55Nq8Pj9eYatKsz97727ufkBAOI5UwKu/LmS90zMypzMdsi9xpGO0tnuA6daWLRF
5PVnoztsyVeOnZ6C/2LnK86CUUlpHSi+CKgs05mPdC0GaA0aiYd35cLkwyKPcDCtUSUQ9aQj2RmE
Jx6Zqk851HEUmDYyw3Tmd2sovrh7mOaTMsSLJ7v0E0W562bZ4TeLNc2fki9ymKgY0NCzaPa+wieY
1nmoX45nhAab0PvThw9wdjJGMZvOE8SQrbgoYLxzeZTwaj2aIEyAPJZn1YvQwWb61PYzqtLDtnyL
jLQGXNWWHBtl4L/Vb7Q6Ojvnbp8+0T28vIX6VpjM5s1WenNC1XSAnEgKiaVpJY/2kalyy58n4PBT
WgeFWGfZW4lAs6v1soyJbXg2A4IhYfqmW14m5qC6OblpATeoFEUYhShtj+E8R15UbaZmXMcqrqkK
YQV+ydp36AoVGWI53wp0vdCanCBhW5BOzVIY3Ldwek5keVJI/9yjlVt7iN03aSvYR4WNqfliB1iO
xPykdqjzhcepYy5lqoEmOTJ7gJodfOKJMzc8ABLWHTquqJ8lz8w3B3FfqRN0m7jIteTnOmlx+I5t
e2SZMvO2G9a21kpDz/Gr+QpZWLQx4tx0M4awZEszPAzZwMDQCgxuoV9I7Jm9RUaRcIqDiD7RWnXq
1/+mv0rIAsi1F4zyOKM86+5UqOcqd3Lg/F5z+GvXM05v0GccIefFcmssSr/bY18992wFmi/oB0Xq
mWPK8AeV5NkrQr9c38OE8p7Wh97HlilPADTtO3ls37NIhm4QAKfEh2rUkcoP8rZXTzGdGO74e38p
zRtS5A35eUTz/Wk3nWnsIHfoB4mQmrrYlYXIBD03N1HAl3uVBSGSZVdetdKVKjK5QV5slrLTKUA+
wkcnO0IyXN7tbuhSfvLfHBMUD40VBcPVPS/fMD7CpTF5epoFg9HfkKLelVuf89oFBZ+sV1xBqP8d
r5tEW+0NjVH0+VeGOXW1p10kSKeCzcGukJJCrKG24hMOjPfoVEYSmjN6ZtBSO3ntQgO9NaKSl+dQ
Mb9+T1qx1/V5nfBr0iOC29bfae9WD0BfLXWAXSqpjGT8ks8pmSfVXVkuEp7uYRYgI271BMxxeLLO
LvkKgRlj0sAqJx99DFh+TijG8J5p/xp3PQiP6g/oqT/hIJ3yqgIb5hnyHPDPevl8XGTyXBaR4TS3
Dqy7AFlyUkYp3Y/Y4wTpN1oT6V+N/q1yEqb7AvVfZj17zX76aSucaKBx7hsjYKDCOPmW0Obde/m/
M+VVilt6TXGuMatSCiZAOqg1Eb1yScUXCeYkXAMCAVgfCfrF0NufGtLQoPnSnWbih2u2sNTnyaVN
13Wiqk8yOOMth2oRtiPgubHjSI2JqyeCQSazGw5oEKX8t4UiIRRkrdzmAeqwU3CjkO+hGVwAE75G
ZPuwIod6FVu059JZdXmHiMSmr9Dp/CDCiBABg8uIW4AIYTPvDQCe0gwyYIEPozi6tAuThdptCw9e
X9j1cStfYcvN4wuigBC0DZOS5mFHYdVcdmifeLvNBmxIb3SogXO+BlgN3lliqH8H6nNOgZ0Oqfat
xok+a0sV+Y0tSCZKeeo9aouvwKCG6srEn+2I0/T/ko0yGnxUJHnMDyv0JZnydrd5opR2ks6qu2o8
LdwtqwghiIBmXfgjQ8vE+q/U+TFkDRBliY4tRfGtbUiKk9BlAdswQdC+vGS5nG/NexnVveVduQ5f
NixkOpLz3ajOjC7q2rB21z2gXBpnzhY7KcSPAibQMb4pH5Kj3QS+QLtas00+Rg0ogxAiQzFccsIX
Yq66tG6l/bXXcHKzVy/pFHqmCjAhv0is0AqfRq0lz8/smSYzoe6cWIKSXEJMGuitVO6MaCCwoo9q
8/jJ+nX93QnP0fiWvBV1T3/QLhko4yp2wc4B650MowMHYI73SZvLFg6WTm7Oop7brnqNaz5V5wJz
BvaN8AytyNml78UyILHfZcd/fnHzcnx4DfmyvhqBg5PYzFjRA6c3nQKUuoi69nA61Jjj5j98wL3H
io3r7hH7GrWp7xrul6ThmBmqNWZujZrO6Miq7b6WDg1Gw0g9FDuKZHg0/x9Oyr22bit8aprZRw3v
qx1eLidIxvDu2YO1cB+d4iJAISkWW7vqBZrz3D1ZWbGW4rVG0Ewab/8XhaYhAF6KQJn6RIJDha/L
8rOl3Mbw2Jp1JDbQdd9xRAgPVPl+Av6WDd7uKhU6MGri0lwhUTAHF88MRqLccJbKEuZQUA8laqhh
mJEiFH7iqHisUQwiZv61x9CEADDPKKZgnPUSg3IjOBRxIok8bQ5nm3UEEee4WxcwDwa/mxmFvph7
NSPThKfBTX3QanVEXZI6FrbINcYr9uz6UlSBOetw1ElGl1Rh99a6iSe4JFQ7BJJE/0MBdTRakVyW
tuUHJMam83TC6pxdoM9fuo0wumHTMaHQN7Sb9FbAbSgFqQEJE/Zp/j+8lRHzpmdDUAfClYXtvMwg
MkhQ/u1l3yslAca1hvAEVmR5u2qX5Vcx3EPdtP6eoaUeF+WjGKfyEjPfhlSPxMLSdI4mAviNWCkI
etzA5k/djEL6BLYxho2pprwXoZc6Xbm3/8GbDjVSEYHhlQ/0+KkbhRdw471k8yD6ETjnzTsThlt6
xOMJAcaUuvRkmdlsyUyxiyaVWSG7c3fCxup6kHViG3/l6cJ1e7x9VPb3+TDR1gv0QaiAQOpFMur/
1xRh97+3hd8IDgs2O1JmqZ64G+JlttXtzshDszIJFs6F2+jD9c+OO7BJ8NARcbqEivoIpO8fTxpA
IyFtxVL7bO7pBCZ6DLobyaLk+PAE4z3TNmX1BoO0LT3me02ev+3xx1GxA9lPum+m36ifcqOZkAkx
/dkFPQMKkQ+uloy0ZdiAciuqiA0kdYaowFxfMO7oubQmvjeKNaB3wYYXVEJzUuidda2DnxsfsBwn
LVr6pEiu6jGlbv8FgK3NGoaY7FCdsiu9WPlTMvwQmOl2PB1L9NeC+TINbY/Xt5DNmG0uC9Eu2ECL
uxbStqNBGptuv2pUsO/3rksGY9HDLvu4A7umQaKb7GW06nzDqbFDrXNTp52W/N900SgD+pE8Wdy0
gq8V+By1gbH5ES0ToVllI+QplZ50AUO6i123AVhVxC7X+6PZgn1A3O7WQqQhFiKBGyd2A2eG3sat
jNXbAYm5lxUyaJybEMHnQKvlGhxSBLayJBbfHtMSUk2bMkZjDiKBa3A3/wm/GJY+U3kcpSSy/QUz
k2HrGii9a+CUfWUNd9HMahT4IemQglOQHs92dtVtbvKkDgTz1ExQ2s/CRK91P+JT8wKKyLPUYBAS
Wnu0Rq8ARe9I0k4V95DATkd0VSIVbznyrobTIAU8OTfcxMrqrvOgRu7UaGMVcGjY1rJKK4TEwVdh
TBbhIce1Rj8NVQQ5oyyJTVn9KU4d7MvpOD3bKMsYtc9Q/TpAu34XF9u4lK8NXMJ9pEivZScJQixe
OTVNbJa0ziC+eeEzbJqGjTvFYaz0WH6nh18oYVSbvCc6J8LURvlYbrzYSvEnzm8NRoVllzwnYelG
LOklNt3rryk0fNrPK4do8sVHfo6ONKTGTeXTSmxKkouZNtpCKxV9Khx29BeWFUo/GcNN4QeIDW7n
TBH25yPzx2EDa4mSYkpyDFBpvTPFIPbNr5Griq+v0xqUy64S3nqb+yhKjbG7xuCnm5A48x5Okbmy
KlC51oN3ajwacbPTEpa3I047lxA2aGFFhTOlLFK/Ki/pe1qZ2jiFpIK2ReK0CcpWv7+eXGWrbzQu
fbhCy/H6NUtn0ztlS+oIQugKKmA+0IZ2wgozRKKB9+GyG2uW794Ux8f2lfcVTf8NzEG+ICnOJyhQ
CikfyO8PorRJgqrZwilvPfSFy/Vk4FOG6NPhstriEtYCWyqKLrrgh/vyjs1GY1urv/WM+RxKfHR/
KOJmynD+NLa1hVQWCzJFN0qYEteyW0YefaTdqWD/AamupuWx5bLpdZMR4iXvSB6eYBY5S5LImBxq
rcN/oHAPMets2SNdv6s8WWYeyeZnI9Zmyj/HmlVWYxuGveym/yZLndpWyp+xSks90kl+1OmT7KV9
kB11rT8TqLJ+zx3HFB0HOfApdc4s0ivIt8fLF7n5TmKMVAM9ZL2EbN1yBKRP+t62Od8bZW5RVimf
E0Br5OWTeuVgOaNfgxNnyVNwRrPR6HudWhH/BJGSx3aBvl5O6PcZFeJN9Pyr4z4xzmYPV3fybAT/
QcqJh5AaErgGA4bm6PPM1i8oBDr5gvUi3rT3apOBfyybsxeY5zZvyJ6LCuxW+yEodRadm6cnDeyv
HPLbj+5uxsng8j3wwoA0wJy1A+ahgkU7rv1bga/r1PGlppCuaOFwREla9+nP01DC74wrgEQCnDlk
ceOuk9/10xGRDGmVDIEodQhwjIa4EKbysvCuxDbYGFabUz8ykvwwv8A4KvdWg9flwJPQvJAOolqM
XRoZRE7xjNRxKBnN38Jxp019Dc2C+WZtuMfYpkYv4CZQDwxBmpgMutwRXeLRsEKJJBdnK/TIyA9W
CH2G8aEJ8CrBrTrDJNWbJrYNGiTWkNh0muQtngvtnaFYXRAJ7O/FH7Usy92YRmC2fRdfD8xbo8sv
Rzlj/W+3RgYDTXAqBqHrzW/HQd94iLGAnLny9u3AUucLC7Nf0V81kBDTMZdqX/trR8YKbD9YQpnw
/+Ecio5xEnbv4J261XDxCQWFmXD3uPWpcN9Kv+8X5Kf7L2uaV3+bzJkIsvJe7JXFxccSx27N8fAn
WnksbIwPor37xTje/ST60tfVDqmiBMr9imUQRRBwkyS12L1i2aBPEJTxAq2tBY3B8lx/lYhvYjYT
v+OKg5OCgr+pTvwT12nfyoGu9UBJ1bi2VU7PIAcJKa6rFrl146Gl/pPdixBcq5b/Cry9GGCjzEfe
pooVK22Ib76lzguJf/NhXv5o/Vjp2NJ7JQeZFzpGBomojOl2prpF8FahGXhc5wKxsQxR1PeKoxJT
Bs+ae4REzkgS1hHBn1SJhexma5eM/UEFZ+T8D1d9/1R9PTLVVWJRuljSajyOTH+yVYbB04+69w7N
0shjkWcZuQtHYWtHlSkHJPUjAPEat7f1UqIARl2Dw7rIyzMDxLN8vBipgLh4HkUfVctJ44TLIroa
+z9M4sekConmbRjQpZLtNtpihl1ZYT+niS0Ws+VQLYmj+SgDH3GVoJb4nbd9JzN9vsf9NWVnsgLX
Uk9F1evbRwuwKkwr4YKkeR+oI4Homc1xAxufAYBTLWTABPAC7IxTDx/MCp9qr3jH7o8IIa8sm9bF
vuFS4Z7QM0GhEK56+c64JQOl2m/6L78gJTsLOuxhkdytAGd3MLSIVqo4wIqkudhbaDkemBVkBJfW
Y51tAxBt0jpumsZe0O8gZZxnWV5wKzfydk/eGiavU9WNZV76/zDfxV9/5oH1A6kidKm7jkzoY3zb
WyycfqGgTrsOX6Xc7iCsyKUCBuJ8Bfj+Q9kJKOmDJeTTyhwoqi4RnUjiLaj9wy0sweQzOPd5hlEs
QOVe9d1b/TSsQns+NzxlicUz1386dd6Yivhh9GUno4WfKknv10WUd3MXrhQu2mqPwDkvKVQY79F3
SGt3JO5nAXKzvJLbO6yww7n7XHf/Bquf6SLuaN6pGTuJGZUU1l66mj5SiMKxEayriMOQGBBfHQXE
3384AObLfnstBm7/AORnaOeRXR/I33+/yFyJRtHr06r+bH2Mh2IeV0WgTARWpMqVSc9+FXgHUDRv
qhCgjAbWk3tRA77YE/Eiy3mhAKkP9S3senP6aO9q8gC/kXVRJuy3X7IHgKM0LIslfBQFrAkAigWp
D2sjxYgZ1Jzjiei1JuJQwPCO0tCwTDomKqiGV4gbOdENPC16InhzYCL36kISw12oAUu9ncFQc9wX
f9R7nM5mIF6E4052ktphodFeRsu/WINICvowtmtHYZ9sM2Ud6rn4xsrpBjUgNjTigBmFrPTSEDGa
yWxUmkWo8gPG5asm89v9muGbalJRA9Ujul1LA1bBvr7LVujd9iYmoc6gdciXj3ytHgW9yMI94lj9
F3L1qMhGIAu20C5fprgUJxEf3APVtep4XPv2Al9H//OQ/Q0GA+92I6VDGrQ2wnk6/YdraCPtCA35
n+h9DX26GZxupftYqFUtyBpy7/hhuOru74GILdDFkv2zkDUFjYjT1MHDul4Hr5TAgrMaVxvc9lF7
i2qk+uNcNZhcWsmskrC5791fzEFOdmWtyzbg4u1VOdSmsX/W8ZKpNEUhvTidTvF00eIHfE9Y5PhT
MUKgabVLzcOweSOOySZDgEQQQ/Ncr8ga47ZyzjnSTvnOWInSK7fn67dS/2bQqYoyyZYuEP5v4S4+
Y+jsTiLtIY2qj+DBoc+19vfWWQ3JT2Wd6/ELWs3R8cGRj2Fo9Y0XhENpZJsgFAx3HWrFvixKZVea
Zz3qQcCbJeiIhy2Nwa+RkPLlwbLOIUZL6paSZfi400+KpDdwzctp5Ctrv5yHZ1IC11XyTlBoTaWE
rF8Ak5wlQLDAz7z8w3di6T+xlA4JokLZRYET1ceDkc2kDXT4MLtyumjUjdgJU47VZIwb3uXfdbyK
0G1Mag1d21UvFLJvMUC0lferXj5pWtG9LO70UoAPJtD6lbcWLr6xFlkQWXSlvwMknzGxA/JuH/F0
DqftkG4z6Z4A6buZ5/TdyVOFrBAmF/cTLB8EfF14nQ5acT+mz7DMoaJbf3+vMevqItw9zgzPnIDj
21OFWndX2Poicl7B4o33PUUNtbOUSzCSmwv8Ywk1SED1xO/PWgDN0NbXCtJpHxMNAvAiyp6/7JYO
71JzXCdNLrqQajszGq9QubvS0WvPxOt62dq1EVD4PSIj9bdxBaA8C+6HKZpcqBnsLbvr19JuN5iX
qCJDHZ+SWHNm8sHHmYoAYasLSQMHncaSTBZj0b0+itSb0DQDIFaj9sVi63FGWZ+152cEcEMDyPXB
5ca6pn7OCwnpVIPUkBKA01RGT3mGu7eNuYtHjWye7IPro8wwhhzvffMDE/6xTUKVfUAdw1+yAVjI
BShc9vqEzYbma3uiqYMIyKklrQ1lCVyTyQ0GNulEBk26TUMf1i+9Ms1e43Thb4lNGvWMpK9m4uBr
c1omkYR6ph0OBKDeuS9SaB36cx3kuHkhCnIE7SSlPaC/gKbcQPx2PQCQjkxXcZn7dSfcEzoc6F8R
OySRxIHvRpcfcRkHBuKolymdcGznsGWGlkhcEzR3dISzTb8sqzCIBc9UOiYgBcsldcAzaOps1iE9
CFsthAh3fUV83YVPK5gR1HJYP6I3fIbKwvqWIIJfN8II750fcE4MOVc7yuhJ/3R8/mS8xBw/8zer
TZ8EeZIF4d++ZfUBkW0g0FRUUvvRWuaEN8mP1aWMa4JGMvDT1rliOMcuVEVuylSO4VocTKUCgMQI
L2XGMriDg2P9UWc0w4zeHwA/e6H07GnVpft/fIuQuHhWFAqwcaF8ezRYrd/kRIv5YUoZyu/hgzpA
A6i5cxbeaUBUFJkz5j+MppqLGMmg217wwLVoHGTbOk9PbDfy/ywVi1tI9mZKE7Cl47+ebkjYwGdH
rpVTniOXYimhX1eO2q7urezKNNBVYyThA6+c0UaS8YQguH8jz+mZtVknbkMcx+Dd2mZr8dq0bdz2
xMkSyqUwOpcLgNfE65lTV3Hd7ucyzeFCsTSRurWNXOM2pT9pKFdWzQ8m7V5CFSu8mYKGyLS/qLS0
Ez7bNKKEP8zGl9E5QER6KCVzfRvlCKYGU0JP5HfTr9Nrr/YTzzdhoUG+dI3d51Yysxn6RJb52VOX
L2aUBzfy7c9S3YMUSvSubPZrcwTK7j1bFEQn6dijRwLR6Hdz/8Fb0vJShn6C8SmXrgqDLRTf1x52
5EQ80ZyHvxkKS6WMxaW6XerSrbQqMQAHjA13FBwezfdJsL2WMCUysRKtZB1kv6+YzVBcg6/y/HPO
T2zi18DiAz8xOaCjVcgl14fUrEVClZaRXV5muW6UWA1aGIUTQEFU+ztPQm47Cj+N5Ty8UriQdZEn
ce2+Ih0HKgMdE7OAlbEwT3pCioj9yROrAo2xmdXrzOVRu5cFZesMr5xCHLFcXmi7hG6Fl/wywTcm
i+s0+7Wx1FY3HxaUuxNSrjyBHenXHnGgQPKbP2qqX6uCwLVaq8DKKQ60G8Qvt/xd+9kF0Hv8x3Ea
alhr56+BiSVNvVnVWTFCmsAgxyGWkkaUUnRQfwNdm9pfONn8oiny7k5a5oHZPvslGhB6xsDanW6f
4+SY4ewVg1FC+13DZIN6HooIS5tnnjU5aMtPG0Wzcy/4svnCQnWp0SwZHKwIppi2FbOpLdidREfp
TsFA4aeeaXP2VrPUJBwcn4S+O5r3X4m5rwc/+Y1UZI7ylr+tKZ9pBUM35S2K1vGK1Cpwk6GVcM1E
IpM4qCejeEDfJiDHGZQgAWXSCZHA9KYuS3twYDBPZY9+sm7sIqt4VVmKD5zdHLQl/j32XU2SKOeX
+vVS2eI8RdpNWK2XGhgUF9nwvW+T9NDIWCZTaVEQNQ8T21REiMAPGHR/+WUSaTh/LDhyKdIq1Ehh
7Bq2PZ7Bc3j1SKV6hcVZuxY/RxA+M7vXuLVgN7+Rw4L7bl3103JFmHdU6wL8FNS9RFul7v+k2VS4
s1R9BA+b++Zc/KiHNLxanT5k6MVG2zLdl12ixfuRqHar568lIpM71Y0aZlyK6IAa/baoM84iaEi2
oBNA5sm+C2ltq14+DSkBgTk7owZ+KheCty4je8VMsYiM7ubU85geF/kUhtoF/gzJM9WXHDVxK7gQ
OVeL5+GvbuMwIWpeBl4Xln1Fq3BOYQ3HE2PELKIVVVI4DzAWwywTdTwOBmw6FlAdT/mD633HXbfZ
15BK7jusNlm++4dKJ5Ui0fpBTQE1GTktQtzrCRIj2V80cGjdprnstmirUS0EpXnFf7aaLmkpa5hO
SBarZThCrEClcTQizC2Od+sqZCjBRpfFdVp8yYoYjTqEkrRWS49xxCp7j4DEQyMXJAXyJ+LvODQD
y0wGcN59evj7CD6C1yNdxTgrGnWaTvsCqCdvrhKbNcrgVYqTPqDQ/wRQspmif2NVnzDP6j6GMITQ
Lmrzrak6LK96zQExMeqgkUO7gyvMnz1cSPCTloWnM2C3Aa7cqF1dU5rb3qD6bTStiIC3RT8tiUaT
esqtw/pbr6iDpwXw4oR9dOfTyxJ+ZOrqsR2+bqdwMttXwhfmoBheIQKeuuhNmUVrLFE9NEsYnZOy
49snx8aUE/pgDeMRUv2CuvY2JVjmZUnHSBP5xEqVj/BA4Ezy3ZWzaUxAhReJkgkMq5CJaP5r8frd
fW0ccYQFtTXVLW+dT3xuD71EdAto14WXBFWZg5eZ4kqkN6XpkEUzgvw8VnwKLGgieW86qpC9cLkd
xM6AZeFkOoofb3hfkzicvz/ThHJgXHfD0xKuQFk+1K51dMGFcN8h/3ZPLjElt/WISuIam57azt7b
cTHmmP1GpUNLB0itaSHVfNkbwn+40qCmPPFh0LXyaVisziRF3HEk2fNhDlAZbISvrqKWmXDIBkXp
qPesVBVz0Uo6Mybt+U9AD+LKTjjZskfQCcwxt6yfXQz2nQyvJdYSgP0xL/dlq4ea6/goO2L4nwAu
NhszbRCSBIfBkEepX5FSuJGL4TWnf3EGxRwr3y1yQRyBYNgKLmNI1fef0O45Y31aBDYFYUNUeDUN
LyzCvMXRjfPc7jIJcz857+/Z9B5lDyBI1xENV+RfsMbonZpxRkvqn0ExuaFNLX0t5IR9Te2e4JC3
HqgPUZ76dkOH7cblBamRafZkskFsoAZWlVuZ5f8R2+O1KUxUfBT/2NZ/F3MQH7V1ikkWOF7yb64w
xnsiJtqfTy8lN+Ka4rYdh6XgbRMEJYBc+RMeAtcXwCsliXGMBH/yMIIV3JyDSHhMsq9zh2SY362u
lfLWv7m0oU4jdZN77n1XgXm2ZFQektM+4zCXszFCP9G0WjQ7T2zDnQeyhj3zmx+QhTtN7MnDfqW2
KI1BNkiV+M0x2o9G4HpP8+5/jHRmu2NyDsojsBj3C8/yDLchcP4W0TpNB5Yn4upZWmHlk/ZQsMox
5ax341attLEfLXxl4z/MULjmOM/yCsWgSytAR8VepYMP/FOcMnTe2xDukWeEz/9i3BaI/pDcNQCL
QlqZvpM2skGTHJnTWsq91520uO/vwgy0A8vZhAROHFB2dYJymFBQEKRQIpzOl9uf/vQO9w6oOb2j
Awd6e3DEIXB5kj/Ise+87tAUJIovtIsg2JJayP81XXf6RYpc6cZSDFVpFGI3SV3MUdj1+sv8I0Sw
sSURBG2MEbiqdsQ8KtlQc1t3Mdjy4WGeHz0pa7VST1IIHgS/PxPpdaVFkZRdMpu2Q2DfycEC0WJU
tjKglK0QQd3jMZGXuDwxZOTp3SI6LunogQ9xS8WOezplidqDW+fMAz95aIkpcNzLSO31HmDeTUMV
bvcRou+3YKFHkmSUS3mSSD0fG4JU4WAR2d70J5GzRnGb9gdk1idOjHxdZoTdySu/U1OPtG6+4ZYR
/AHMWXjkORDU7CBgtDNtikpzTi2lEmamtINWTorTVCU3oVZVMMPLX77TB1OLPZeow2M2W3YKTzes
awnbbaTjiczr2dosERh6WwLQ4igFaJnvfYAq7yfu2xmwgQB681TOKOcr7zZjhnWC7NNUU27DEXam
4wdlFzn/BdbBQ9R5pK7bH3uETsrQTQv+Z4jh4hSdwwBhvxfBFE4WX63weLEvq6eoFqbbpfEfQxWd
gcYbaa7ny3fVTmL+jgzWyyp752qWSBWAbEpLDIOfM8owj9PEvE/fLlbnhVrxSq61pADKzSSRs5Io
ScQf1fMMwrdHp1hki41qnM7oSWKuL4YxhiWJgdo4rcda+Pw0jYGJfkV2KDn7HEQZVPEYeAiUS1iW
cIEDON+DxU1PtYuCEkPEI4xzwYg7Vin9GkZU7FRlHQF2RBFh1MfI7ZST0b8hfEbeBEjI7PY7xzKn
N6TymIzxbdQawP65frOXEnpiZUyKdQ9cQR6UkWdRZkkk8TZYjPaQqLemDK2bWv8P/9Ng1nbF5q7G
59oXXwZvGzzLIXsWJPu/hpqzd1P6CZTmH8ASBMNq6p62LNYs6N/0urJwTl6wIKXhExvQ+xGE3X+K
hpUckpH1XyvBrhn4UfOn/4kCZktvhihSRvmJ/3Eb9o5meFZ5Ig1H8uVOM5koRSRy9YD6Y6rD+3FA
Nt9RwQ1iEivmf2OfI+UuQuRHnP/JBKockM34rniF4W7Fa8K6qTUTznJaQAHOGDN2WYx8yUBqs2Zp
6X06OFdVvO35iabbRm9KnJbhibGsZe5BZmIivzL1/eK59S6IrZgbgKqW3KNhY8IoPPZuMmmzY590
Msrexp9iSs74mrbdejxthIYvq5f6KVapKUZqw/AVpuhKIOanpjY5S0bqGM6RpL7aINzbcoc1ht5T
9t7TO82dZLozr70rHcc4SRhR7iBmtiaGHUIJk9Zc8D/GBuauAsN1EayHFYzOxA6GP25QAKG22g22
6PYRLmVocqsH3MOPBnpkmB7Z9PZ+AdmVoQ4V/kVKZlLq4M1dlVW4o1mr1uNcrNi55UihDF4CBDbi
sKENqC9iKJTKKMEv0IIR7tJ/nuJwVewvTyLa4DGy+v7FiEfK+bBNrHyIQZEzfKLTvhZngYe1mqdb
kFs85UiWHSnGnA7UUh24nQ4wXZEUN5QSP+bObG9PCSczAAHk+SaT/sw+8SU+qtF1ywkmYDoIBBz2
vPbegpeLduBIxAa2/YCqPUGPqhvLKAfGLzdG4em92UwuFRcoTJn78srQGELdYGZUn8VZU4d4hYuR
+XSwcxNueTx++gD0iBCHvSXScgsh25dk22uiH6vdHLyz0Cq4VGQMQ53vUN+VWijelVi4+ru5cbNZ
f2sdfzpjAbhDQZ5wgYGOU1fjfqrf4vrczey/mrmy/3kRDJqKP6HzwUK0y+qENm+wFFtj+A3RlHcu
JVO4A+NT4ffCrUjyP8az1srsLi9fq31NlMwF7igvw1hc2tVllP7BMDM+aE19oFLRXTmDLsmqoUrv
U6iTmzgsrHRdcIZbqcfjlTk+vyuNS1M0MtiJJe7rLhxUHZfUvcc4/naNGElGkTMt5zonMujjcowJ
6jLoDvv3ty8VxUt3s7XvyjLxpSJQ9K1adlDto+gsIRazIBJIcincTwPGoqNC6Gv1Ncy4jflp5y0I
W3POrPt8XRttkr9LapIIv5/gtpOXiOH0JEg6j9m958q/Bnms39NEEE/mY1/MciKbNDuATXWjNSdo
hC6FnDqs+BMLxGwimlTOEEJmFdoQzaMC0l/gyq3eZncRWdAdJoZh6nq0HWJvjlagoWTAH3QwobgD
+kM7XvSHPGyQqv+DhYaCAl3cpkHw7Av7qjY4i2uiZvccT1sEqLVp/qjYrEyJXA8KhCpiAnRjjdk9
pHQqVWIRw+DrX18lx+PQN1tcEOZANamU9XwCdnSIKSm4mAOtNc4IAqzlCJthwGpveRMqo5Oysfxt
fl3/+fJ3aAR26PdZeyquhGXgaZRGnwCHOHdDsrMk6ShKhhwds1z75sZLKKwFt/PsGkxIMgdsv8/c
5YydPHa9Px8v4jLy7njiX6ITMQ1J2uFF67AYR5rjBKrul1q8s/Tt3Mi/JlQeBbi0OzjtHRwyGYus
Bm7j917jkHIJk1Kg7fzH5HKCB1w5/XkFb3KaPnXVvNpCGmazo0EqvTtbx9ZsCJCDWFtGNgEoGooJ
vp/y2rLHCjT7qpJQmJAh8cQaDcJdv2ZAmG/TOPoIcdZ1tfDeG1FapRAAPBHShKLXzMpovvzkgvnk
K7DOc6y0EOixQABMTKt2ZfEZwUApcBgk7aH+F+NJkM1saKW2zC5ZcFdYX2LgQjDix/NGY9Am4gqm
a7ARVJxb2YTRfplOKmaTrhfSo/77nTW2Mt9Mngir05aaiUBISyA0BwhZl2nr/2qxkwmx8/vR9+5i
BpPO3eE2kPN83Nv9al8c1oPnZHH+Qs9mrIHOWVhOmPqObZJy1hJkTKTLcX7Mo9wRUREzRga1cytM
M7+S/EI4xv7F66MQnScV3fecpV4arwxLPL3yO+Rc7e5dFlXO8XBAoxqn0sf7jMSKS/GMudPluYcO
/1TmRVps5o4p5kFZfQmhbzaA9KQeE6OVbecbfikw6v2XnNrt7/h6erUEHuurZpw5LxjP9lOkmIhC
sq2tH47DtQaaRtfs8jnTCIjAV8bjPaRMHciNNCpWx3DzY7uti60KqHg8NG2xKSfGv7D9VLmsXdZq
D0wKkW0fFLNYlkH2S5wd1IYzxlP83h1wdm/sXVYM5k3NcR1HuTyNuPUkQJXqjZ/2sgGeinEcoogO
lVUt0+BkzzemS6wXqabWMkEhF0pBBRxlcs78THQwDEzykVv8caoi4mhb5e0bpSL4R4+hP8z85vg0
9FHohA+2d2gx6fBPTCez3EAuinQFlgZ/TO+DpbPNBPkFcWg9HSC3CJAA3svkzlRxpHpaAztwb71S
ZMzvScIlXFRRqsrpYvJvU6ZchIrKYgVxcO4VF/cfOByGj4RIr7JDAtuYt1QdTCGqUR/B9drjkQDx
bxwrFM//pF49ugvrnG2PCaHJkkyvPq4TkCA1PA/HD+NUSOTsWqMOjOaJyOJmeTaUOreJFIkmN5ql
WbmwnpTx6ctKSg6y9JBzqpKBeIHKgO2MCEHL5yUiZoF9glkj5rA9l6xBgBumFEMz75qLiH1z6HfR
n297ry9M/1ayQdYq/TLBT9yFxYpZMsejKvrxidrAg7tA4yOO6o4GqAUNWA0xytf7y7Ano2yvKIN4
NsZz0to8RnRqSXXbZNwR2UwGJdjXb4qhDJnqGgx0C4X/zruuDYYnT5L3dJHWNS10Cm4q59jJ8NKz
m67iuKc10owNvj0EqWl4j/dEB6uJJDMaKOexq/Jnq/z5UfkEXYImqWgqVTXMffiSMJNE8+u1xktE
ty2kBMjnZbVgRvXAr95gb06AbDk0T2uBVYAH/7nVZuKmY88plwbHABsqPTpbHWxq5ddmNXhv/usd
+mQmTXYgBsfb27fo4ZOTcq2cWsi9ht4vUw7GQwocDeFloNTnuYmqqd0OUOvJrhITxXdXhBcQzMks
BBc/pc8iTJZy8RYha94Q45puVNmiHtcBUGGmpe1jTzqCC8koOm9jDnSSKgsPVJEVJ2HKMVzsa89q
z1x/tyIfEIeyVtts1RBPnTbgeune+HJL4uUxSCPC9I2lYS1VlRDhaurllJfbDAoO1WcYU8Tm4B6x
Em7BCRUzs+wTDD25lhbzNfxU7cjx66wnEW9u5UVzlhN1r3vU6V8JcfUetgqA/TmqP6n+FW/pjSks
9xpua7GXohsDV6947jqEi29ICKRv3GpE6Cr179rklypFkhWNUrTJHyyipC9YgxA6mGFXAUDmZ3DV
6fycyd5KZytscvZt1nK2dGDf6TWCIiD0THw5eHmL8c3Mju365/4XdrekfBqgM+mEoK1ff7We2WUP
ats7qimKjC4tshSfvZKJfqkrC257aQZ/hM64xBtkZhOSUq879tKN3gB2ssewzNbtHC3Dd5+KlGd9
jAUt2KP/dUl/Vv4TYdkG80m1hQmHXylYnZwuxKV+2bFOjrdatUA1N4NXTjk0YD3SqPQiwaA+vyxz
KNLQO6Xn68/xjKlfIrB+axanQ3nO5ZabOkH8Kh1UmfEjAa/VhH4hrrmaENoizRc3+QTGd3ouKmRf
azufYfkx/HiYMH8ZFW4831whtJCuzbUu4iy6nGELgjq1KWWo1jH5a2FAlvhDiZQ7yQEU48E20a+o
P8X2raEHMDDEezpAxAdFQI/HQUxolY9yuWZQsNVXKD/V01/qFjYl5gNWNxzllqErWRTiQ1ZOWOzI
vCDs8o5DSs9/GyrOtWm3qcNclI5/f/43tiiymTajUqRZHnFcu7WAyPBExcFB04W482nzeereqxI2
kjovWpvWXHx+EHyT48hmn3l4UHE6lOu26yZeIpmTLkZMEoDi2eJqnR4GiXIayhvOG7dKRQC2QUDb
2GetekdzbE2QGcEbdwxK5wm9qmWc6o4jTQgS1YcePqD8sy+OSdBNhfO9rvkXuLJXDhsZ64+LfHQ9
Fmrq3EYk2tHi/696pq6X0LMfJqkgCJFiffHrDmOcTlO0h2tIK3rjTIVLSNCUNEwZgtNu1eSizyzU
fBJCVPqDeB9Aks0b2/d4Hc1+Goyd4iin8/C19PRuwZ6rRhcL2b8pEdoEBwBtdlxAlT+yxVsfGZwO
AVIza16sDTGIt3XcVKx0/oOrkdx9Rhys+IUYjpqwjLWC/lkTkkIqcVttjGRLt9w1Vb8Wkab78a/O
arpoDxBqwwDMW25Spmj/LSVzCnOsMaK4d9oZZZUVi7niTe9fES3sB9LW+BgmU7tmuzpb/4rRtuhk
diSFHAQ35rtoBb1hN3pogQYKvKH1tHVfKpdoMFSp3v4QQ/6WqWb6Y5tOF2jac9rnnCQdEq3ZpA4G
TwVJZV4CbgmKbC+Uhe6Zo9p7YoX09p+Y+tpkuvCc13IPIekuE+iF6XhMf9XKnHnYFNxNLYKIYUiY
+RXfpjN9YluDh7u9VbiBX2W4xOCjazG5adYdnvGOA1paGCVHgFKXdtP4u/MnpKGGbmprymGtI6Hl
YRmFSUJjPwm73PThwmkIZ0IvfUKtRRxo+MCHza9kK2RRRM2bpWDrpwMF/5jLf2Gsqtbil8mCa6pW
W1j3mHUm4kJmEEpQq9otlAb9BOq2UF8qWMeFnMz11Fs9+A4MfYVaHunb1ziXJjhz6U2VnRAislTZ
TRHk+fc5ZVUKKXF6xtdg5E79lbaOtUAIvD4I945nO5hpSSKapqmmgHXxmgoSPEYO5Ok+S+JITIqL
scvFhypChoOVg/roSboGgPiz/k1BgzVSs0+OPR5mcrpDdwZgeH6wWKncJIz3UDrr8dmkqW4pZLG2
UMndKciCHE/aqgR3A+xcR6uEu2xSSq0ECwWGMmKWGl0HmRVu9v5+bC9olJt3pHA0DTi469dgNJow
O6lwq4TEecCb2DVMpcTVw9E3PTLhko2unsGC1GexTRs4DM4OCx/GHoPc2obiNevfjNfeCX3fadTR
9Btruact0BAqe5JR9v0Bsx8MUGASmgXheGkw6OqNVlJ3ZHCg6PtWCZKqIaWuI8inmE8fQbLM3dNa
57TfHAwGDmbZA3O0xPpu5+2whnuQ8tBnzR86HzYK1/NrNF6fcCrKCsqihWC8r0KEiFs1BL6J8tcO
avauITpiV7sYjB+gkPve+YIBSzkY1uPHPS7m84WE/mTndHqwui2jcowgJ2D7tPbLKe3NW3Rrbkmh
oswb5jwoeya8235qeQB5J8I675S6YAlZTmTFav0QWMLn219RoGs5J9BewDtpuhrDKeSIUk6vdb7B
C+rnHd7xGnERtNxcxhOXzZrSNV2xwJ7lRmRiUU1QcAoTCHj6VMwmH57D2tuVvRCeeFNb3pufHmoH
0hvRujBGyLEwPE1c39wHUpAeqiDux0i0uKPbUkaHwB5cBrtFRUY9cBDYof0Iq4PEjp8PMYjQ3Gyt
QrRMgIGuMOKR/i6BENqbnarDF3iKHldfmPGyH6YBl8SOfCy/gCx8uYX5yWj+2VdKPivDoRAQGtIp
ZCU77ur+q71qczkx+MgXh+8zckSQg9lE1HTy1WS+2Z2k72MQI/tpty8mcftYTvfzAg5d9SOb3F63
j5DGpjRzUon7BePCnHejjD83JdkRr/lqi7HTFtp6D0eNBVejP633buC16d4ZxrYGTpDEZiwuvv6h
JAT9nSd1KTlm4ktDkd2D2qts/w4RMau2TOrn7zFIWzYF1wgPKT08lfler3fdOQOOOVRC12Vlr+Oi
mF+Mpj+MDtWGGXhMkWP9WFTLf3sC5v62KTtpnFSb9FG0FJkoGU8k2Jb2oAhAiK8TxXJYmnJyFAgg
YK4T7FLiBwYqJzzfo1pf0rmaeAUD3gIjlgXbagVNIqrXGcomgw09JVOYy4uddpQ84R2MMn8VdmuO
OXp5hxNCCy+yClVeNE+NsmOQM+0CVbS7R9CRUAwlRNJC7koEUDvl3sa/pxgnUFgkWoXj/ay/IxNJ
2Kuu9VO4ktHvKk/yCmvZcawL8ofNHulddejIWwMtRrNA/VT+KACWoGmggoAwzTwLLxkxr8mnVmpg
bvQFyxSrgHRDuZGbBorHcg65v354LsOZLBV41/iCF4ZV0chVs1g7Do1/Fe86YCsaydi7UwT0Yfhw
E7L0MT01TS42pWKAPaC5Jx9wmFP6zLFxaSsLvRT4qPcaYhIgUlgX9zSMcCnsKYJ6gi+koEgCBcEy
jRVI9+QhVqCM+eyiXOAnjdH2eQIKU6FHRTP5mIMTjgWWIGeLQcKFaMRtSOPBW7C4FUC7tbpuHgdX
SAi7hQMpnH+rgSn1eWwB+lVO99owzYxGvpIpyyLt2YR1IFZFA/Z64gYLRzFGtUL+VlVktpNqHDVE
FN2JLSzIdPf8l0b8yqbT3Im8lCAo7wy/R6bz9JJRqerqF+6RCIBtNYEZzFwW3uc+DHmQi0KzI2GL
0twyUzk9dHRTca0WceZzbRPp5iecPiQNsLHJFIFOFEpLLeWjv5VYHrJE5CA+QqxmGGBvmcAWNWIi
20t8V4cwr1tyVPybz+zCNU8NoqKLuqIjU4r+KAXxQytbj+eKCeCNpufr9b77o6Nbukk8j5INjCEt
UeInUZ0nHGsbkh0BMJYLF7zW/fy9T+pz2EfHtJnkMcmYy7q/EEpP2x2R3D2mgwg2f0FaxXQaFDho
q1vCfV94ptzYLnZTbJgY6967e9SobNCZTMOrwyzl8nJQbeYbXnzHqpCs3yhZaeTAQ1S+E3UODk+X
7bwhJ3LeFu+cZJLxk7T5HmrKEYJRhW6qwqXKErAX9dHEMYRPrYqQRtanrFlXsTLWCtwKjKJPhTlL
3fYVJW0jv6/pGYj03MiA3wzefz3v5LmotV7FD7DVS1U/V/DYku2lI1yTbdLm77+WGobbhTulPc6P
FLtseNfcxMN27FPl51ZpreQkNpVB4wPAMvzPO5dRUR4IfdUO/iC8jzWFKZ4V7xnwau39P23fOj9L
+H/9PjJAjc8pTLTpKupebo2vx2nQncO5EiKwdeliUE3aFLgjKuDQEb3D2Np1rBspYlOjacpxXSkA
mTfoVzMxd+Or0kEnMwmeKLPg081oNRWw5oxExZYaqMDbepbIsUGmeupv9a9fTNi5JF8KFvJP9Jd+
bRfNj90JzYX7rgrqKq2IkxpcHNv+kO/0uEVD6fc77KhCnKT0OIkPz804HcxO7O2C6JFk57zcTS7K
i8/V8i/yX3tj7JGUFIR3nidfvU3MUkO97TGcmrqz2zOs7xiAinHfFnIbA2enOceUlhHkamflC5sv
XNG3dW+pTjY6eIVgRqDXtIlU/n/qZtAfo49oC/s3I6RFyMtFJiDK4zozTgrKKR8ZSlsS4Oek2koG
9YxBEV3onX7W958kDhTaNSIIpBeJe1aFBAbMH9UaLFsWZ3p1JtU0px7gYtQnRV72Bv6CTYIjqInS
Nqn2DBD870AJFwj/FU2Lmgh72D2WwtDkw94wYiSu/ckGWsaR8gXi3KKpRoUwsHk8J3mkRD2sEc4d
l4K+OKl4WtcDFs/KRiGbrVxBSFyy1nvx4/oLIzsnca2nhjT31bwTf5tLWRN+8IwSszhNowAXC5OR
UcZYEYAZdLhhwaURfpjkaaEA1X0sTPVbsw/I1kjri2/R2JA0J+TCo2Qv0nb/jtVOu9NkMHd/Pzrr
q45ZW7fC+XdI7etczYN9ym74HCizAYlQgfKttvLodxv5Hoscm2xpqDLeaOg4b7F3SCtmMqQAKFJo
uEblVPSS2Pm7rt50FoK85qwlO+UqIel4dz54N86w7c9wJV1PAX9EX6pIp9d/Fs43tPbm7MK4khr8
9N5YUnJYgGWq56dBP5zogbvGSh4emPDRWX1lA9GJJVy+sSy1hB5jF9qChkNKEh3QOrIUvy4YdNA1
nwUACP6PzhB7siduRhrNWNjXs35Iil8kuBCqBvi1xQMrKzRauH3cr3+5iQ6qYmANrNfw9ctTNK50
xh8NSjAvHcG80m5xXnOdhSxAPd32vt2Kidw4aBKuEd6UsWeyOOmKe7OCWBAQsZDA51RHG18ifHUT
q9CyGGY+wzL4cnxv3IVcYUV9RJb74WNAsuAJe4hbVvLg3FuA0UPfeHg1pZdMSzWEsbvNB4yDeREU
BkO1ztC7+BIcwdCvtTfAt/+YeUvvL4Chy2Up2/p3DVAKSzpczmCTl46yT7+ngehOkxwl9CWUDLwH
fTMcxwOcgdIFak6CO9VqrKmF+QFMtRrUQEXBIyyUeeA1SAOQl8LbIoBPSf5ddtVE15KZB6qBwZ+i
7IWy67HM2w1vg8UqgiErCDQe1ERBzgPrp3X1wSt2mTuliOgrGCeYL6y25+zfBE0aT4uN1LMzlK5o
PZQ+yOddpv9JofBhZ28cf9f+aNoup1iODnyICcyGVKh9GhWgZn6aLS91yV2Z5vd4clRpJIpudLLP
bUcBrmJdPnhgPGxTbFsDHGMbBchiw95qrVK8ApD7ezuGXQTgDJP4zUWdGd0ns6ViicP7iDNSDvax
ANYMRGo6FT39+t8T/a7/77nRK7j0jXwHBf1oz2vdqGYRF1Okonzmtf/ytUSzajENXnm+AnpV0f8e
Zdfz64czZcbSjO+dgdruv0pR1XNvlNlPzeNAEQtTbu+wHy/enmv01E14Pub4O6yymjvWfb956CSb
o4ZbrDv9acrqhr4LxvDpbb0VjC3WyZQJhUNRy8RoNpQCeYTv4VvCtHlL6VDoVsjMUCh9FGzT6O0X
BjhjGprVvADJ9BaS1oRccARqfik15NdKfILeyJIuwWy3Re26g3Z2AeYDv3Prw7eE59IkqHd0F0ZR
TKbSmNVHf4q+7HwKOmsKWxODxK6xgsW25LI37fBz482pP/btzWpZ2Yot5KM5wjFz2eNl6bGD0t3e
7aeZf7E2ggFwz73BGbE4oRHOBYXMEAvplrOoYMjGIBcbars90705Qjp9UKwaltcuVSBYs5bImA4E
9jBcw5TxkK3n3gJV6iUooabeI8FF2CJyeZf2juVzuvyGoYN6QQCfUJ/ii+qx4j2nODnv6TxVqgQ6
8xm5c6OVYDlNWHPuokRzkZoV1ow2FzOVlkse3pdbWpL50lOILC76sCnOcX14o4HT2IwAVWjrM+d8
Y4VWG9cti04W+95lQBxlB9OswaZ6bJQ2QbuECcmD+mqCiZQ9K2Lu6hGa1N3ncEldAD5MdldVgaOn
w40dguZ0f4ln7gqMemtePhuAA27mih/ftVaasKVtVpdUxlTtUQ2dwjflv2ScIX4S4FCaTFJhL4tI
hyS+gtEHt8yQVcD3j/nYxjN1oID7APK4b/Yl2YoGmJmdwYi+XC+/D7kWYvuEAG6xFwBgI/gSMVM0
YbbZvULM6IKt8RBH0BRrxVxWf0+dZIztLHnfLnfWt4taQp4dnqhF/Jo21moUSWUH2Wa2SWZj6zRZ
dD3geYTb8gwuZpT5Zeu6biOWgCiS68AoRmO1y7KBoLByJ/pXlHvHzV3fGAY4A3ms/E9pUOxKfoIQ
5iZsPI1pl1muPSiRsY/nfJ4HYS8d3wO+fjvGoZv6mNtgLftGox0pUajIRIb8JS/kuVO8mj4z8Y9Z
Iofk2j+DLvGoys7FyCnh/mqbmifRCBwf23lM8xoK1xHw4pZBsiQGXMgeJa9UURIyJPSG7v+bM7N4
1V6z8A7b/EP3FMzV36YTpsALgtGcXzVFNOBgyRINLK6q7jPv0eXLocEHSTjpu9xcVcuU8MYbnM95
l3quyv78xHAHjw00jJMf4BEooeXOr+0anlEgSXa63EK2itYsKvYEEkhj4IT4pvjscgJiHS21or3t
H29MO2LB9M+EdArVSw79pumwke6NwdceUi4mAmaV6kxDx8N9iup+3+n8qYt7Cca679jVZt91UpWu
EnTJW1p8PAo2eZd4pUJUBikEuPbgJwo7AQ3kP8vBjbHwo13po9fmvTRHyjImCYWANk+MTPWg6bDV
eTja5vSm7Y7d4TYcY/aoq6KxxqYCr6vnL1fwZb6K0IpNQtC++C0MCz5/B5ZG3ElebLuqjG04gW13
lxSmwXqzMifyB/BfZQEDT2Q6p3T8U+YDyZNYPofD1ywXhrfZCGZi3PnoClQkKS2nV9Nu0e8DUpjz
v6QPUQaPZOkqNBWHSBYEuY/99qnlAEq0/N3m92EKnij+AWMGBsIdwn7ifYh6hSNAY/CaG/xd7t7q
KiP9aRuMFVWgIuhP39acjF06EkrLNnEZT+tshwIMlqY9WVjtm4Sme0WcqjmMG4YZRyRIPCXzMj9T
rS9EPvksvClYfvxPT1mRG43PMaazsnK3MkqHFcNbTMtFrFOY0/8qcBCp431ZYGoBZhktQYUe3k4z
NzFyASMiSyd9eJdd8r9XBRW7HOB+lMBBIRLitwAEUO63f+bBqMFV9pbWHHBqw080zLR5+c2ol3qc
oYxuKVy47miDiVNLGP3Mw3vbXotizAMdbTdYuwV27gka2p3QcvQU+9GsOE6FpatyZpettCdfuDH+
Ytr/cAqE9sbhuw50Z1ctf+0tjIuO4FOliue8A2uBe4RU5TiUPR9+Xoy8WYIWskXnH6hMiW7Iu8eF
sCCSmifQlo8ot2idtinCgwyJV3xHebCNpNE/RhpYXRjGp1jzQXMAnYR1Ymz+zxCD7FBhW3rzZSBR
FY+mW7q5xSi2Wioyh6KtqEN1N8nputk9FVhYbmf/iTXgdxVFV74ZE8vmKRYruIm6AQ7+nh/9knpd
j3Jqi2IH89kncWUF8JOnnm2YUsxyKvg4XD/4REIv8PKQD4RCbN6XmiUdJH2x8AQhKZWPwPU8M+me
xbBs+yLPPYfDi2OEWS4qvpCh9OgtLOcJ3hbVQwCzhWPq51OrHw3kuvNgd6kjsQ5B4oI/Z0YiTPp0
hEJXUdfOEDS6QmHi1sngolieG3T/KhFNAr8rccRhKWKMYa09uGYXrxE3/TsNvvIPVw5F2FEec2I1
v+T9Yc96smZ8us8CWxirLQfDtq4mYtbwHScxuRdTYIBJDeDvpWpX8qCdqjVQoKqpwFbvxmKYZgiD
AWKV/n2Y1EjGrJe2gj0tn7+NW0nxYemEZDmMv6LEi2Vq8XUhK452gKoNQLUZRSCd7rb1/AmOwHhn
D0//JhSvwQmu1qqBcQM4h7Yma39jYReD7EcUABSO1sSPubyihm9SnYnt4rp98o+wT0LlbxXCut5m
Csuxj6WpfogBeqHu0/slE3wTibZCqjWa3JE2JKJBqutN6UWUtIRvJPd15aimaKdqGTR1C11Lebtg
Xxbf7z+RrtLNF+Q2+JtwbXWPBjMDzDWTksLYVfdU1JQxVSzPOX+tZi6kNCYncLrvmZrIJrKYZOHI
34aF9sHcOIkpGwu8c6Z3ntpJh9+9cOY4KiGFQbJKziQAK/Gt+ey4sARj0jvlNtDZJEGK+ioQ0UnO
rSIjyjiTliiStYQtmbGBXK6Vo4yRvhj1Nta51scHLWykncSbFJ8wCmdXuUOaVPh6Xmw0oDTgFZZa
eHRRZWPKmsn2kTLqOSntj3JyPPfXO/86Jx4S5EnFAjHOsEC2OpqM2zE8TKnkIpwHgG8slOLEW4QD
LU6V887ZbgYlhAVAinuXLA2PiOqbfEKsT+sP5Ym8p9CPNKtPCbrnz0ebVUAbopsB6NFT56AMWZ+U
+MGb/Ms661mrgvBHsvFgJ/fQ/2Y8qNv9yU8nkdCpKq35sbamazmVFwBwe7mQODWUQa5jTNAI/Nlc
XuRSP4Zom6dpC6h7QXkQSXMhA+v/1kSDt2mRe7Yf+pLVLX+MB2niIde75hSUFrymsrZ4ki0sZtZC
2X2BNNlCxNxr3M+3aRSAAQHSR4aWPGh9SF/hr9Mj3zkCnsRsJnQQHfySQA3Z2thEac0ahepX8w1I
bgzIN/k8ypxD8Ma/m6yYTyIS113Y6/T8OzTg48AaMZFtXiP+enb5XNO4LPw6ZG9ahFs1zw/AGSlO
+TPKK7wqcth+ScE9X/3uBOrgwLAeYq+IwhWltT4bZa+BN/0UIM16gTIBafV8EjQ6ltb6r/AG4GM0
Zrf71N9EcIHDKhxOga0chTfZ5u96WDoDNockq63kLHOubES67eu31gDl/MSP2kYRb7F4/21uU11W
mNNuRvfjoZjYpko2hCy1R9IvrBLGxx+AH1B34yjNOwB9ecx0VuabRhVPbEV9cW/VhzYRkGXwnq3R
7ycVDzgieRS/Bv8FSO2R0vPlaYOelL/eru6adppoz4FLiNBYiCX/gTa/8bkwd5yaFP6IMY9JF3nd
8iV6diqI+G3e1eH15PYWgNWtkn2VLp8BqNmTBCYX6DnFThM020yRTolrODqxv3V9Q4Id3EaFwNBB
hBeq839hojrUk1nd1UpvWk54ZXFjGh84Z/6f71oy2A0qPhQud7b5eO46F2/Ts0GjQiYPNkK8NxOi
sLm9Mb6j8V6osBsDZVHa9jtk/JpgWft+XrM4T2SPpKboNSsMzgPbrAfK9c7i5gY0unNrA/PxeuLn
4e8Ljuz04gXWOwd49REYrh7MgQSOodhMchawbAb6i15+X0xItPjD2tUDhcWT/mbfBduTPYjVlAG9
gulqlf31uvPIhLOmvOAK2hdXA/ZdJqpLcDiIcM0jH5tcXJtZq79sxSbL8TifzNp080BU/mIyhqW8
lp1uEOtrL6PKU5cGOqQNMHO/hs1uYY3YKN/D+hjDB2BM1okkLvgsrQzTUJ1md7Nwwi+VXT4MOWBY
vIj8po8nxph1Nwny7mOxReSjnpydV2VwhUP7pMcmEgxGdP+UYytbDSy0+0yq1SU5qoK4QfUF1Ei5
xMScXwT80KcQH6RdGzPQWCkaP6yT5EXoaVqqhgaYPWsGFMgKx1N5IEQag/fkCrrCKHZV+93aMrqM
qCJ9+rirw9Zb6v28qVG0388bg/+Yh6iwJwkIvgQSAozGOwGEwcXs+47gI2jLHK/jdsKJ1rGXF5fD
rhhohh8SkvSgDnE573SrdRXzRp5cby9FKNmfaBD9VslCLHOojfHyu/O9slnYJ/TWcN5ECGb9UwqR
T7p7r+uItiNoAMSgH0QWAM3BgVkaTsD2FCWkDQFOGpbn+rs+ruTL5jUHgyS3uSWv5/7kLOFQMgsY
QZ66yl8RgZgBBevX0o5lTMnMwavW42L1sbB0accXZJuZm7zel8xQRfamTBY4qA1eIUZLm00KyHIs
CB83SWlCA7HB6xxlCfUEZYSNWqVUfHBUO9Fk4yXTLTbG+UpavZ9WYXNn1ta0aY9jQ4G7sqBi/wBb
jlDtSi5lbVjm6CFR+YWDNgtZLiXIu7rP/mz04K2mLnNAXD+82uppo7rmRrEHNn4FJ0GlfF/gZb6s
N+KdfJdipJiKLMoTWALKjbzjuwswIdfZF9PEWIrRkOsuINoPyQbGyGb9cT5D1n8WWXswY/3zE6uw
v8/HQ/tYHTtdtyDQUXXRHbN57z2KQhTcONP5K2H5lFgEYPM41TgN7XCzE/m2kmg8eApm7HSGAWPc
U2raPzbe/fl0X+wR+G82Wlq6ZHHSdxWOGsv4gpBz79B8SzjcUt62Wg/nM3jeWTg7QvHhDDdOhXbi
4yK7ftx1bXGGKE06qY+TJXZD+dy15op/czZFpenXVmmR2wLbKvEIQc63HknGwQy/Aaj270tulXaM
LFUOJDno9WrUJ+21yykJ/3Pz+WOeBwl6AHgHkeQrcHdZx8O2xpXeJ8V5jboKPPW2UxCIUSPSY1G+
UppIjWvygwLJJ0LmvehtA3rIJgarPr1KHNdtYO1XrGX9b3z41eLhZQ1chXnbU4nfgKPWiVUCgxYB
ZUO12I51T0hkGqn9OJdjH7ZjNWWhaOOcK97kS3ZXCI1QKfH8nliulfcaNMHosR0VnOB6+zDjeKG4
7biFeLLoTTw6kcxB/IA4myOmMKtFXmEKMiHy/zNC65/YJVUNGwE+BjmMejQaPCxDuOD8BBGXz1AY
XmtKnZGNncqGUJEAw5YRq0kPu6nSD8Vj+bv/OlaeVcKY9His9YaHKz5rbbbLxFB+oKYI5vS3b2xs
j8etbC1SAUc7IagCRQ+heqWTj+l6EXLJnxvaag+q36y1WpGptBdkIHotVC2aU4ypaJzD/9hbjnLi
v0DlUVQbcPq2WL6iqOBWGVUNHRv8pjrCMCMd3NaUZ4lkDYKySpBWTkj99GqXqvMGnDl6WQIP6QcS
g0/IqI+kkTKffOdXTviMW+CnwYzUbgLFth9npboMa/KXeDtGn5nm+jP37I+1lSsSGrdKlF3JWtXQ
NwjTQlfimuvpb4Ezbr9qrbHBup5VHmSJZSGuwqgWnXqd7y39EWizoinrhbUmsXnPABpSyZI3Ygz1
UyoT74xAfMqWhxrW7BTiQnTztf9iBjQKZEwUe/XK19mnbe53L9wG2SoTwiDgf5Qv8h58buha+u3g
GLWWdurKdhBQA/0nz7AG0z4suDiKmPhDHIKdwe1FV7ddDhMlO5CGt/KaIUOxV2tYNpx1PGomId7Z
uXCaQS+san5wA2fZTyLzg/d9/gmtXjZS6L65y/ITxj0NowScrErVIEpUXQgmVC2ThK0+05q5D6Du
Gr7Qvvdu+EMZxLL07uDnL4ktNu6SbhRCiuPGqcbZeQyVaHFPp+ycfq3slj2DJjM/vjw7b53bdX2F
NFychuSksp+I05zHId5i+S0YcaxufX6L+8LwH/ELm+Lmfbva+GJ2zQ2899vc1oPscHr0J8Or0D9X
i33GxXB2WXL7TVKllAOu2YW9NwahNcQu2ZUay8u88wgY3akCYyTnfX61KEhRq1bXtnQmVn/eYrY+
/38Gi3VrLWY1SHlAvdUfOgUuOodrpldjfa8ZQ0+exDIgEB0IWcL2yc7631UlQSKboWcckqIHrxUR
il4ikBor/SfgjmLghEbS6e65rHckgwhDB5hh7FK14slkWUnQ1ztHNXxAIKM4CLmyW02/hKtkI6VT
G4QfdwB8QOF+E7OsN0NangNOD/QJEZ2YQdU9yuVnC5Tq8/Jg0qMhoD/asIz06AFYonz1O0GJRcZ+
yyyigZpBcKPuTZTiOYgsi67h+2JGcWS/Yzz2k6iEIa7FcWmG8mHT0LoOu8WXaD91briU6dIEQX5Z
1qkXTPMtz+BTmyH3SYNNz88vph+EmUy4BlWGwxbAMMgEd12oj8uhMAVLGrZ/J5Di9r5CMAx2ySOs
mIJibeCOS5Hn1mDH4EOizAlLHRzY2NYLJpoTRuFrIxWCNUjVsh3O4RSpaS3JPRCQmFWZcmHpABUx
hfV1+lWwiZQrCwoAL6KLhrKqzhV765cyP7fC+gOhKhbNRZXeftet/wWCxYXi8tHHikQckaFfhF34
HEIQEJnX3N4V1lAtf6NgB8lEi7QYIQWLzv1gTjthpVoct4INpd3ymW5a0N9QLDQRvbyGdUNX/BlI
vr2vW6x5cz7d8hV2MpOR+xvVnL/q6YIIKepqZmoTAvBw2lln0Hey/Npv/Ayt+CrfAKUEgmfhzKXk
wJcZnFQ+EDRIOEVZA05X/rINha5o6wLoWwtz7lnILkwIgJ7IwKF0b9Kbvk3estwywlkN1m20gjXN
ufVfpjfQtE4rZLJH0dGDqgiSajofX0dHl9J8ergiF3X354eNxvLzHikquGje8xsMfJoPyGRa4ijM
0SrpDH0rO7E6oplkIBZbUEXZl9gdJBcpvzp34dVno1x3NrBYCFxzBAxpgYaGggJ3sZc6a73ApfVn
BDONJqQyEiulVyCBV5j7H2R7+GfP/8IwNpzUcei8iY3OlS8Kt3V2q7RA6MvHns7pK35VDfLl4kU1
l+EzMTBk6sROc9JzVr++YdoikzrwVQ984XdEVWjFeSega0IxwZlnzgtFz/KHhGZc0dcedq1HJ/vF
lFLER4NIfy1mWtwMOiC+2t0dBrkezGxWM3BQZs7nEoso9Y+qKFhpqLs2imeilvrIZz1M7C5y2T5B
JuWziI4MgYBOarrVFaNsp9pTLASXFEquyHyARWvOYT4T+1NM08RYKcubQ9R7XwxTzJrj2nwRiIIn
iu39dDB0BEmVtUq95UnVF05SJpC4RjJNYfhwQX2naXTVnQmwVui1W6hgqZtpvipqCzE8mH6LjYVu
Om7+mDby4Q63UbHP9wiz7yJSJq+UbfF2l3jr6FfGj4rhTxCdoD/OIdlDGAZH3pXTNuaGizz0J6XB
Pl5z/D2n7wB0cHLRStovXr6D48osCDxpbHb4/r/A08YimRAg2idTcatby8TCWbZcC/YyQpScB85E
Yjy4Sag8fWbcdwT0rDkv49sTmXbNlPgVZyuJwkOcIzp5sELjaq54u9CHbge4Cbs0AgCGgJWvx/3F
B5ENb9MkTR52L8+NF6bCX56AWWlkPfyMKRtGoZaRpndvar6vonF0W+sk8uwCPyTgcgvkWHk6vEOh
Ie061zhf/EEM45AKymNsjxD4rabR0YjpaQYw53qmabYimPZDDZ7ButJWM+wE5vqbxUxLM/GteekM
TiSVDW08rN1vxNQglm2ikitcx+Lzri1u8GzgIFPhXPzLzMe6Cf3Gkk8uO3Oq8BB8Vf6LWZ7yclI+
2UHj4N4xV2UYUKj1NH8heUgoJVBg2VM82XqFvh1+9DC5ho8yI4w9bgg6ebXXYcz6aarjeCy9SETg
YFPxwTkv6Epy3CEfrmagKIHpa+dRhLxDPnyCSLiBhLFCqbGSxIaKYayQmAQ7qLRfs4OHhRL3lHyD
RLMads70opUv10odXaS2at0qVGjhOWHorNxWqYxujuTMBGNqgYkOf2uQacb6lkOjp6PCF3+L/FuB
PJ9Go+h9/KOyFTDH8ZSimuTL8Gn9K2TdnKrgzdvgFCeBwCpNrvoAaEeY56kx3eDE0fbBVoNVvUPM
L0jDr+M6kPcWMn//GU2V6i/Ys/Tfm9VQ2IFloEtRnh633O3VDkZZN/XcWQEL6x+JZJBDujSxnWmJ
xS3NghELVPROxlMY5gHhO7F6607vm42ktZ1gBvk4NuXL0I/wAmRMRB4pNbM1EL0rulntZZgnziO2
IVd8O4tI7jG3DiPp7tB3ZDOtvKjhcxX0rKMLmc+im3GsctWZgznKYWK+x9UzKi743lK+EREvR3ux
UT3R2vaMQdzhvhPFy+57IL1JJr3idqahHMjK88Cbb19enCuU9l4TB/zhuqyziM2gu8UG0QmWIknj
LHh/qGS47VRi4bwvnTOLgDPsCpC5UYWlwpWhpzlzZaeOSsnaoZwKzV6hUUYoKbWiPSrOvvBJ37gM
rcHSMbJecFSHdqvh0A6Kwd81jcPmOTUB4aSEDPo9G6xO2thjsugQRO2dKUDXxAXLmXePL9hNsTGn
nIEEFKJxBZcCGnM5RwHCftZGwlBK2VgSsWn4+7qDViUwu45jwO345q0kfZoKwPpNuplTklEJ0vJP
Hsr/dIzy4KIILI260JI4XguyniUmf9tChvcKuoPBAdIhO8VlUfS9ZxRV+rMk0sdyJzSS6kDTEQsy
SwM1TMzeSSXU9rXIIGoioLL9ANT0JTkWnARQ23WEFnm7wvU54Y+bN+OfWERt9/jGzxBgVo0UpbJ7
9OiX5UcwA8J9wPWghM8CLTUzg/gTs9fkZWo9DUm3UmbWPeF1SKxRunKvhWMbGwpTDcwhe3vs+pKW
q8ivdWpky3rR079cEd6QraLxMQx81bnRovorQGhOkBeZpapAyAOEdRPz8wNfI7l4X/ZCXIc0Tjg2
mNsV1ZhjDuIsS+URBxZWcP5yo5arSSQT0XgvzAv4bDRi1z3lgok1ck12Tvml11ZtmXjlZGwiVkj3
loHhwDJpe4H3+RN2PyqeAv2hWAIFi/79FwVhA9TZXOzkHUBAOXMiNDncubp+2IyqLMbU2LB8RDF3
O4QIjuoLWxSx+o+VOqT6uhlWKxxlx7rMr6kZHqMr+M5ZruCZDmJaosxhPcIEmjgBchfXACNHgYOv
kWqJ9D+FPyqkfjImQxRqIN16xz6nPjyyFdlnscsqOtib0eBIIvWNhphznQ3vxi0XMVLhz11rmhsB
hYIuVj6PeCuycMM1cNDKLsNt4QERReRaWGJDgn3oChjFLTW5DYGH4L6/E/59ELWfW6IAXxCj4Jz/
cTMh2hd8rRIxQMmiKXG1PAdUknihIqKhTVsMZy6crVivW2W841oqjJuGUvOoyKYCorSIRL9xiZrL
IFYVhWP2Me3NmIqc/2wNkn+tAqSaZI97c6q3Uyq/I4vvuv03Y+5mcutsKskzCm47ERwKhs1smkKS
1j2ohWcS6YnDEtdnfUjoK4Y0v4IaP31keNCVqk878Ng517WDIgg+GBjT4j11aQ72bA9IqqbeAKVg
z5AIMlBOccsIIb9Cr15TwJGookaB2qTTOEREaBkG8X4WVi92BRFpTdx1TFIHC+o+kLCvXVT+UV5w
OnpARUV8c5oehJgQcR1PRzW+Iqo4TATh286W6a6L/W/6Q3otScoBNuECk72KlkTK7VVFVkR0wHRV
O5BS3amfeiSRQZwsLW4i7/NWxSdE+B0PtSAQbN4TbCfBh2kHGkLAp3eCOoTpZlTF3gRfw+Od4B7g
Vp/6MtcMpp8ZxXcFbbxdMhvtnVzf1xIb5MkRg3ebHlDFiWwsLoZH2wj7Ng2AFyVIDmSYspEwgjy6
L3dICWGXNqgsMueZNbXxyiIR2yFH76ZNA66LHDoVqnd/Fj+AJUe/yYpFp0mvhRcc260tLjzKQskW
PLqnOOIdSXd0oLbFi8tBw02+8dLjZrz8mIU2JgETHzM2OzWNEh2BOmOvO7xnHP02Xsp3lg40+bvH
SGkw6pZxNy8exXgMytu3R9FTyzR2cwA7BAt3w08nOUYUQY7GcMzqoU2D6Px5nkE2QTf3Key7FaVO
DXLRj2wDOPvcUzYPfwPhEpieuOvvJGDjPFgQA8PC05j4Df7Uc+sXs5QfKhwSJhy4TzDo6oJqPyju
BYc9wak1VWrA1CajC6wKzHsQ5PcqeZifHYdhbXr7f3b9Vaayg8wZswbUeyhMKYvHy5zGFK9W0G74
gi7tNO/UjmlHqsM7aPM4CLOprHhNmDWNl8MEIMG1VJIIAWEP/usxEavhLC4m/47Lxjt9vWCVFciH
wNLMdbqPAA+25Avt7OVUDy2x9NRW3BPaSMpdmzCUF2dalSTM9ZChhEcC8dSty0o1HnCz/ih8Bop6
lHHaBFJ9KlzhmOFbYfiKtlBZpPOPayaHqML9lF1+ksxtrDs8JFHALxjia94eWNMgbj4rTm3WEPjC
4aE5fEPeXcwHTXssvn5weGnow2Ys5cSH9mg6tIIzar1cj+wn5BKpi84KSAwSe7Pw2eBT+FCIdgHk
4rkKwKDwXn3ETWhdpkOmJEIJsSst6zvr4t2IArYoOG2o/Rx4TLoAAdp4NPMlLrBF+CdD9rG4WICf
vd14bT4U0zsP1EFfBkp5zZJOPjy5NbcgY0Laim1NB7UzgMqaUr/y5gkh5ypx0UJmMhB0tPNLUAS1
NJXxqgPEPfzwzYpAb8zGaCe10cPx9lGzvH8ylGsaY0YCMrmIiJoE9PeW35jHXRJBY6enf/zCAqIL
fSQQIe3nSUxlZKF1UOHJbp60UNVcM8VjxXJ9sBrDjoWuWIVThI/Cu9+FIhLKkFaynnP3A34aM4ML
a4/NTY+wX0h6ScXjwneZVObYGm/gi9Ko16KB821aCohpm0XFW+XYfAZLzC1zESUw2GWbXH3BzmGM
7dRHQrmC+88c5SyIvZL8QlR5azRe11BQNOqURfW/+JLYpJZ53uoDJC/jVjQgmLvGvvVRgzjBfpfV
Buas0Lu+UFphrLj51bBEbBbbx/1wEBUwles6MzVYOMZ7PCmq5qz8j2Agoxs5KoIolyou8TTcDNVE
1N/gl8UwBX2Wwh0sv6GA1OscrkX3HKW7VtTVlTnS0S1Vvz4Vsd8Oo+UULf8+k2o+nNpVF4SscrvD
xN+jh/L/TDoNJBApOklVaGQ+8UToAXuYWO2VboELltnm0jjVzHRxfkn/g9Sqn6PZ19e7HoXCzjrC
/5Sqzkr6D5EO+Xcm6rkR9FuH646eP+CmhOxlU5fW3lwoI+e1KwbOfOLfDTmsXyTb9qc3dmY8zFCJ
onMKtWvffyCtNmpV5CbKTJskNZzaqSmwwSVH+YLDwR9qDIlvvAwkXh2j1tH8ezbj2qdPVPizJlcM
LJ5hJRCBfKKDiME6zfiiYH3NDnrinMKZmby3YtlSHLDGjwSr59gL+oA8Xha1CrHtxgLCNcHkYe7f
5BWiOXPe+szWQH5yedU7NeDoxj/fB08uxdeZ6kVBOiLmmD3mZhOGdCswTA9V8TQh7+Lcsvey7hmj
aGHW4SnJkRrC5+11SZkS+a0hjrdRG19W2Pu4gnSr/nGb5KMqPy7nRCjPBt+2ccDlFHib2CgxvUr7
kjaqR63yu0zTRb6RrW7r4L5EDr9ldyiLj8qij1rkeARq2uBHxaZnTnxSXI4EWL8Z34eBwzSCmqvW
iT1jXDd1NJfKZlylqCaVOjyba0zxEcVT5iG/wMwJQ4oUvJXTqDTe8ohByYuL2bi8++mKuSwNVcVD
n/YN5Dy8xxf7etrjd11sUscBChq63WuMBhrXyb2ygQQonOswtucEeFb4lhCvELGXUJNbTIpsvJYv
X+/jq+pVqAkaIFrvfBdWyeq5w43WqFITRTfQJEdA2vjn7juUlQQeSLh0iJ6d/bp5oJ995FSjimqo
yXdkWqxnA7s5ZrXxfra9ZFK26MfrGb4AP3sa16HtvBVjzR1CJNM5Qse8e6dAv2rTRMj+uemV8rBk
aFCCr0hQxArSg2h7FpzTvji98O7sww8bUkHJ95ieOHBRj2iurHz25A6zPbP+09Lu5oYlIiMra1kH
RnTVNqDBlGKbDXrzF3sZZyR002I3JrIScx9kZXTxDNhCpKgljZbVAy4/k1VdCLY2PE6S6KbTWjsU
G5zrN9ckXM+ISDjRq7l189r8JngUTQb1y5rn/mxLc0BTCJPR0Y3MDwp1f8bSxJu1VHAl21LeQrv2
kklRVqUInJ2gGPdv3B/8CfeBSyY8ugc3DbTOVOHCfONAtTjK3M2Lf7wmowg9yAePwsZAGJW7WbQy
L8+cfG8WjJYhDqTk0eQVa+O23i+04nzgaEWZ0CfPuPTfcYT10r4YYs9+PiEz1W41CC3IeYoF7LuK
zDoJtoYUZPC8lCueyUZ+g8gAahofUdJHP1WPyhJHKO+uU/h9ofevQXmBQS5tj2KIiTdXRppza4Kl
KyygC+ppnqPyJvVsQ3DLlFlL5VQ6wkOPHHtN66SB+h6o5pQhfpYLf3cwhD8JcWy2Dd5MAjqpeGVh
HITxRCBgwIaqC+S8Lz8kr60/aBsilYZF/cc5imC7JgS1hqhQnmNrTqE+73hVWV91r/dJj2S0nDNx
U1+yw+d7OscpxrQOFwoGYiVhhAqMjjd9Q2e9PrYPPml+3Wcd/YDWyKxTnCR8PjDsUKG1E5mg9pCg
ARyzYa+4RiJMD+PGk718LkOdsygXIloP9tGS5iYV7j4YUtj0mq1jE1zI+lw5KaMxebZv4kehUtfG
ZOH2MlwE9MFVTuu2j7iW4U5XEZPRRy5auuRM4DZWtx8ul8RzeAH7NOXjRDaW9wMj0d0nX3NL1S64
lxSi70Qz7m6k0Z1WFHd4QdVxZt1irZKUuvujHuni1ELVQ+RvHl1CVuMXAvTz3YJcT3STSLcBWwwd
/NglrjI5nwqidXJB0GrTr8QtV/U6MMRwlDUSwuWVDnIufYITWuc8RR5OQjDbxjB0PnOR6Q3pcPPr
Iy+vztCUyQiVhDG8vjUsiL0/tkA2esgo9nuS5vauywWkG+nz/WqiiLDtF2HjgU4WH6eJI+jcP48O
t4vugyvNju0gn35ZjY6rp+Err4AawwD7vDYCI1oE7tz4yeJqK/rGwf/Q71h4m0OQFWi3tYK8hMzl
8fWEXbSIz6NZbdJ1ogD9gv/a+38ZO1P9Yb4nqEZ9ma3QaQ9QLg3VP3X0ZMz9d7ZziwSBN1aGAC/q
PAbtjK1J4FRc+Um4e1XINgGJRWKOKKSlxKqgDQ2ux3aaknN1Y1Th0M3M4GzOJtZrJv16efCcK/F3
6khjKDI4P2OlqvqwOEs3FzM8qm/lsObME86rTkBtSEpHJGuWP6OXFnWe3uESLu2uWF5AIAxr9yia
AdwnMiXm1EVnP0Pr7zbZUXuwe4N7izjor9vJYwy6XZJa5+yzV0QUu7i1RXXb/wjDBVau6F/MvAm8
pRE3h3bce/jDGjASRWBA8byhv+LmtMxOGzrVzZoiUJdKAxjTJfA29KawDaBxUA3CMsilKbjeNcV4
TsYj22FpYvNPgrlr1Ozq7KQLERhtzvrse1ksFevTb/uTMCK6jK1GsNlldURIryHOj2n3CYoipz3V
Sg5vQ+geQnGMgY0zMatI+tMatxkbd/fJMRbY2dwHLZqWEMXfXazHaRs4R3Sx1QPgpueaeiSlSjnY
sq4YtvZabK9PTCMbe462eK9ngUuILovQExaMy5Ngso9mq0Aa3DCHoGtB9Se/UnpH8XykqhE6W8l8
NMaG7/K2Is9Hp765V/LX5C36uccT8jozkmCOZcSYvH/mTSwPsoEl5N+AdcQGQocIM5SFiNKowaYw
oCW83FkjVfTiob0KpBzIb4KY1vIQY3upoCAvoC50tKX4hiJDZ3Eju8zj2qNOPGm16IsBmisBimAA
VWIApSVYBPtw2i/PCop8oJXc4rOLN/lUj1lXzFCPHibQG9BXi+K8J6nO+n6/SjPFXiFfQO9aVf4/
uPTxOSeNe66GLoSRTRANCKYNZOYOomyql1LNPVzSnXGq1sUe95/umRlho3n1CMsOkCaKCyBMMgWJ
QgDy0IpZ2wGKVjUix+jHZrO52mzZCxInoJqgt/7waiHZ4OCXIWEIdMIkB+oRy3F8lGilM2SnvOl+
EdIPHJjjVkaJEOatoyTgYoTUrHQpi3zV/W3njOBOCFegztX4aG7abhEBgJe7/JxlBlF1hgO2tOFI
JIPu6K6czeTEDiEedZJkCa4bQmh53mW+96rztkHUmXXRa00jnInXHmlC3xMyviKdoZWhemV+1l+Y
G244rRVU5xoDf91Hbsxam/c+LCnNELb9aaHino6QzLuKH5hdI82DFzR1WFyytAowH3SuWBv5sk88
oq2x+tjrU4tnHA0KekTiqbs6fqJJq0+1v7PD/LoLawq1K97JIpQSvT3UhuXAqkgI1IOUFub2zu9U
gMWPqopaupBmySNcLYaW0QTT1p67giKQG1n7LBjkKSMm3sP5f3yYm06NXkOF8IImWDhtXCtXtic6
jVLCNL/PtwUGhLvbG5p7aCrj5rtkyeq2kLyX7QN7FoNWuK2ywyq7P4/zvrE8B30sRXPMi313acZr
+q4ackkGcE0Tespe472F68Brp7yQly4BmHcRp8qmctbjFdn0lYFI8kzN3nLMNPuvj1IZyDfGdUfN
X39Y8/Wtfu4JD5DXjDQJ1ICqlH+csMLIGhJbfTqZCy84He4g90GTrqa+5kEIiIIfRXCG7en5wXf9
ld7d3ufEFh9X3T9qHmhwU/zCBUYhevJV6yctkQCG6GcBgD88RWH2YFS0SvbQnPECcpJzgfW0u6KX
hkqHDfFF2EFZ1i1QCNnogK7NydryCiMOt6FIaKuOUc2i167t0tJgt+3DFJPS0E9yv3Bzy1URME6H
2lDY/Q+nbm3kShZeEQcQRD3mM5o08yiTwhCCh1YXl2qbps1xqRuWVFrOTXtzQiapSN97wtwt3slJ
oSIMnSeDuH11kYPrjJLgwM14UEpY3ErWf5CY5KYj1rBckDu9yLnaKvYKB/hn+eJmHsrekq2ewPsh
e9WYd5TasqG7c1thvRisBeMv7Z8AGvioMRbwYU+JIFKP2+hj4ZHlg6SvvTt9n1G1IANuqI/joz5X
pR0NdvX2HPpJg8I9fczTpzPyNW/3dN45a/VTeUZTKGPXsBqkBplTaTJA8T0i1bKnw0vsLK4ptTXM
fvYcSJBflCvJFL9teOUQ16+8Yw5MqDqXon74x8GStmN302dQ7ro5JpHFyqa+sl3QnWYZMfHh4MRU
BVT4+pdQbIn/1XxbpzmhnR/0bpBlbF6ltis+iJYGMqJ/iBngWhHL4EAuX8rXZGVQpPrMWpk1R93s
be9UEMv2dB0e48A2+LlmAUkkfWos7CP7nlchamKJPaYVhT8qitOx3aXCNb0Tjrw3J93mo+eFdx6r
TzI9t67GEyu8fi9yOqijYS3qmg2pWaE+LpBXLwj7AI+rpVF0IlP0gTQBUyXCDlHQXDqJpWHAGJxg
PmMJZL+JqjPz9htIrUUQJiTnqH0LtE+Tp201E+txFE/TJ8C15bKz1TXDEP8yeddkravkxqcOS04m
Z7XAE/XDCmLCjl1a/mHTwnykYwLM9+gDWosk/X3cx8mJ/p7PiFr5yBVf+PaU1mNqeozhWYLNNhQx
9M1WmQUfMHEBeAzZ7W5xaWOCzJSBi/kLjAAHBG/mtL70vtSKyeTmd+9ogex0/jSIm4yhhA6UAXz4
u6SSdfFhk9tBGn+fMosuMQ0bDqFpQC9Z2qsg3XYaxSCY2Pb8qi6dibsV4d8GO8w+wP+D9y7AfxI1
m4Qu/YR69luq3x9osIeTo/tk2a0E1zMMjFvkZaCfpdeco7CkG36BA4Eo7KTN7r3tg459qTF2xqPA
TfbvoOc7hI10o0eHhEmKmGd20Z5IVnAysz9gFsXuZFBhJujCWjCk/I/6cIFUUWUvfGx/7aWB8e/6
IpRq/OE7Yz91b0HnD7eACnmvmiFLSkqJg8BysBksFPzx/LWl0aZkzcvjiqknpcw4quDENg/1R3bv
beBMWENDdR3KGdsybj9d+5CFFrQtmXsnl2hG0hOHfBWfc9b7rZTB92sgrRKF3l/vtvYu3JfyRqHj
aaYWwAnBZAKdCGgNeTWRTDOCyrXgS1Q3Cle//5n3KOBgEF90+wyuQJxTt/VmQPEWyvW8wNjak2QX
FmjpJsACjb5WPC2IUlUI03fDdvbdUUefvNwIktd38H6lp4+4mO9J5eGUjkI0mmeszqUD78/2WeTN
AppaVK7dIDr+cnHYb7/4FmCHugNQHP/5FCppXvzAhLFjKS2QombNCq+yU5ZU3+hYY5ctzSbSGlBY
A047dfZ03Rv1VWG5Cw+P3eqGb2ET2f9pNW4TC3XhvSRrI9jFAfGdK0qncqk6CqZ6gtvn9SNUv7mD
2Dq1VJ2/ggGNmCofXYE3TrYb7RWCzwmS+Ea1EdXsoJmGmnK+/3va3BhVr1M6nWbidq0NquRnSxHQ
QXiPRa1PbuZEDBfKG/Omp84jOK33COt0M6YhDiML211DQnGr09mv7CJM+BwSudNDmBu93kVI+DYz
pNMfQz40otRvbq8kKlfuSnrAvi2UXOGHCo4udWdJP7OpSkBhc7EBb61Aladlxx92kdF/r4O2ukjw
jpnSmZyR/eaSSDi2BX8J8MUUbaBY0FdjaQkFn1+4yNIxcbiQqxY38b+nkZg9l/u7fJPR2fUlRX0J
vd5kL7iSSJuLDG5IB71dVPWQLy4wxRrr9QklQ6nEh1Ih0JwwVom0vBG45Wh6SO53PWv0AbuQYdkS
DwBapr9vxxIv8xdaKoqaHXAmtKOg4SOSJUbuuRfSyBnWnhjVqcEfhDyL0Bwq2GXTbJ1h8FNKDl8O
IWBntxR2XpxBIVNxd6zCSwJ4DydxrMCTTN7Eh7cHcXL/0g6+4yWez6ENqi5MD9QJvwc2xk59k5jQ
zAViEQw5hb4rDiPQrIfTLCuqQwtbPisFKCVmhGxBexV9/7LjsIbKVm/3wD5HV2ZI/cMtAUYZxylN
jbs6UCb0RwFEyNGQIzjiHi273/srIYPE1ulIy0s6tOCNQzc7Ysm8NXx3d7iJUazMu4Pk2WYe+6R7
ypPrBL1o/PbulgqkMBNQAP1qDM7q3UumiT+9xyzy+4dxq1XeFVn/Dj4i8aPRsUpCN2Qv3UGCawa+
TnIXjAbimPB9WTrGFASdvtVekVfOSrCkR6rbvx2OaKw/sis/t3BktqlXwKh/kiR6vd0GF+l5I3/Z
GEG85GW4knyWmPr0vCEHwlZlOP5TyKPW7eK8hltGcxJlqtPFkuX0vVXDsGU/taZXz+jEC94/+Jnt
W50TF7nri1S5W/lfk7XpCrVrvv2ETaLg6sz6BSO2cSVQDubKqqVUdk6Bd6upNEsHQHpzDtQjUMCH
cIx30rk+B8xjc69zU4H+ezVcOVUV1btcR9DwR6fNo5Hes7ra+mlWWhraAA/IisUqrPtDvHmJXQs7
3QwrHvJkPNlh6yvhFcm40PlpLVcvafoI+Cn77hNFoyaQrtcxTwYwCOvelsCqLvVnhbowb0zx4gkl
YapqghOUEPo3St73gnFqE4n2+eMYE7/NG9N5eQ5Ya3aOUxSQQW7TcpYHOdCTsHT44wMIKSg9yxOK
AV6zgjeAJ4EGWMyhHZyn8z6dEXa7UYkztcklW8LswlJTAaiQ/lhHlb6+xqphZjEYciEX56gYdan4
M8qColf4vKXXlI83eEvQsXhgITdCzNKQewOv+Z311T0LciaKiQjv2NaxX3mAwXi6jk4Qi3/2YYID
mUCQfCKx1Tqd6k0wIkAJQLArcRHYh4xGme8O6iX5wHi9DEvmgeAus2fKHeIHpakVXj+2H/8RPZTn
64JkyJULXS8DJs/DHBtQfAbWck/U0mG5Wo/UMegtEt6btIH+TuA8HFZJBCPMNjY7hWLZQ1gCJWwt
uGZjTUk9pNHKMVECm7wb2h1zRMA2PWIfbH4Uhil9b7/a0yR1AEvKoHsZwLdTat7LTA0zletxa1Dd
pQ48TjIiQWTKv+Qt4gtnEJJgk+90Wt1amN8CNosOKPFbHn51e3UIRB3kmU7hkQMI8dgkao6PrL4l
HxqifaKFualtHvdfUmhD5wEhxMu6O04rHRDgyW1qMp/hITX8MAIwA+CTKpt+8RAEZyNkrk8Jc+Wc
FRAiciwxghXBzR1nfNygE8Yr7E3sZZRc5v1wXf3qq/3Zl7p7mpt5mUzgo9aDjCUcK3XBLwnqEAPb
/rsim4TKcCX5BsJu1CPu9OM/3/WsR2dj3mnfiguwzJnpMyF8xG5iFM2V7MnzQPjcwufAEt9kJanZ
X/6j7Reg4C0Tl+ZPWeJoS5Ubh8X88K8Bp6ksDHYul34mTYBbxKVnPRs9IOm4u+fuX9vl+OWfpuFV
OdwSEKPcr9pPn7/LkYa0rX1rhvASQIloGF0zCtaPEQTyzJVF39/Rfs3/Cm0nM8/bSGPHrxXPBA5X
PegYxqnk/h0XKc1Ue0VY686zv+vcaEOYLuGY1fEymAt5W1SpxWIGndO88M4OflT9LYU5wonS5DHi
lcY5T9zDsOhy7HW9rcpulv3gcZFVuGAgnBEXc8zfoxgUCAKqBxhDL712dhM0li5U8CPzQEs6yq0y
nJ9y1rDkY11E7kOI9E27kkDINgP8rLV7J1pWq4B1X2sMmVvDBstmY0n/okhJJ4lBlDvpCE3iM7T4
B8HqJlTEk16Ee2VZjsd8sRc4NkiGp2wpRuBzE8NSXLXDxkZ9ve7CUVUtixQAzRhOt7x7qkjMsEq5
Wi0H+NfYU2Rvk92VWgENe5wQ97Vsa9hfHv175UtZay22S/LcRamWxiSQle4I496ayB8LQffWFket
Q6j5tlitraKxVMP5QTU7ynQyJRlUs1xLUMcKVnqqLyN6VoSZ3hO5dOUc1XYCENmqvrH/PFgq9lWX
QhdztUzVdDPYqtvLyOaA5qvymMTU+VEg4u77ReVGGTdQMq//AVcBzmcy76JrJZBRr142Kb566IFD
xgdDsFjX+J8FPHPNHH/3vX1ptW1/6YLkwxbEHXsAFnKuu1oZS/rr+EiKVhvmqM4sPIRIU6ueybmf
cglUSlFHZt2Ftjceiu4mHR/Porvl5n31Z/gbK4RNHRQLi3srooT/h4F7q+hvMDHSFpH43LuwOa6L
n/oHRFHsAy5kbbu3SgNMgHG88E0WFSvA7FCYJ/lO3fHyC3cOQt0ZazCBdNn8Wh8VjMg8Wwk40yx0
Rc89GL79L2CO6VCKFb+Ov/O7Z/AzuZJX8IjcPASlsPsVSBFhwyXx5Zdu4pnJdcr5oXrKRF+yBrRB
2jqM2Lp/lFyVa5UXJB26tlkZRE/fvMTlX6wU8wey4D244AURgtQwE5n9ujWkcnUGOmLZyZ0IMNYb
1vL+Tp8cYcdIgIsWseNu+v8QEO5OypSAEv0p1d+S9d03bHINBFYsbt+plEY+qeikdiSwBcaLPe6e
xiEKsWswV3n0QfOA5xWPlICwifEW269Rt0yAF1OU355Kc1FF5fiLAubsm/qox8+wNZlcgg/5KpN3
UNVhLV2Glu2DPcGy+d2Q/Hd1AWK2bk1zXvQyhQLzr1U5FPJGQ4k6zEzy/mk4DhnWqQHV+za0UHW5
/Ogf3AI3toLB2RQIPLB0gjnqlQciOs9e1aY4lbDzQfn3mk2unNprsdfqK4JEBTa7it58Euz8kuWv
wIsdJJWAQ4Ln4ThZZ1kl12vvFFLolebOwDNnS10xbF1i0+6+YKcijEq3qVB2UjL+1kw/F8Ts5sLJ
TgOSp/WhxLjUcig0CY2MRDXj3J7/iGy4IPzRrL/RP6C2vrJhJmZcObcuRG28F9UOY8MydfB4gig4
XCqCsEdXYpGLvimCDrEGgBqp4WobosXvCGU5o/CvVGcgqL5aSh4aPZobLQi0hAmATLpz9GgOYCP9
dnft3TNoF9zQqe6psWq5wDgTFE2I2TFvZhcEQPJF0iRt5pWrsFgQ12pal+/r9AuCG91zh5dhTh7q
+tA9Hkq+/p7Wipxz0wVGU3PXLX4ZvGYXzh6HVdt6Ks2driM7ehVG30ZNQMnv5vxmM1wD4C4proaA
ZrFrVktn9I0RZuc7XX44ErPcQCWba9VEUkinkXSqavfgILApiZezWApTX815dRaSfjxRlrOGctPT
MXCVrAOcgYybeEZpVIyApm0PAiouuwgvcC8kzS6W1mFu562pFoiUDHCekxTpQ5FYV9Lva+m+NJyd
URnKm6gjOiz0FRnS10x12A7cvSOglp+ApEMZdGNcQrR2VfE/MCKb4jukXkiCK2P7JUegIpWsqEut
YHtFRAMZokwqciN5UtNUy5guyG732Zoq+ANTBiJjSTp6M4eKiTfcqex3dAuibYHziTw8J2JfoFOB
CsHT1Ul+nJqlJtkdEx5KZBUEx+p0yyGuO8uw9St+40MYhiCbXw9yMlOnQeoDUkguKM8eljKFmBKW
UoGWpVZ+7Oc9nSg8c2t+1vaLG7VTKnE3IWgEyy9HdfOJxROF152FoeznoBIDdkS9R1IUKB58t+cc
Mp5qFC/biEcS6jpVMJ8e97uc+TXpMj5iLcisyBktwId9kUe1D+fkWIO6p1FGLZAQHrnJJbqR2pYD
MuZlZrI621pzvn0ZHzGIkF1U9KdyJBJNhaa9tLv6Bee7nfmZSnmk6/KXbsZUVwdmyNRQmybgvwt+
NbRgloLrjkLIi36VwzDSRfbC5KmM75mSpu58f08AU9CQs9KvRtidGT44cK+/mwgg4DvELMXi4/XJ
0GC0z+uPrb+07T+PjtBwZ5+oYROENoRwipoee4t2oVZMAOwBzMdYvWOb7UDTN0AE4JowmhTGiZZm
m4Ud7I1kKVB7mlbE3ic8zsEOctBQjROqoSHm4a1teGwj386tNYxWPg5DyfzUbTlveAd9frjrF7Us
4htVUAjtJEE2k/JIKj9/ZEzPuSVDW6kC49aHeMu5PMJAW/UFzFwXVobKW8GHV3Up+J6eeOi9UWjY
MVahkUHEZzHXVh1g+sD72JV7vJ1GGe1QFiJF/txnpYQpk6p10ZCiPV623ZPaQErPJfpe0uu54Ldq
0Zo2sf/E/sGpByZzvYdocImDus4PrP6hXLqDP/WozHtPz5io8E4cuB5cRvT4hgwlzxFAY0usB1/I
hUsFjhcti6xjp9FWCQnleACfwEMjpt9M9pV6Mi0AuZHJVfc1DlSwBajVaTP7X8GGooykmORlRTqx
Eyjca3ROmsxkAIU9MlrCK0oN9ou/zYUXomU3baaDJDBwROuTDuCOb9n5hC7AuQFkgbCXsif49FYm
lNBCgPbjfF8DdHCbqV/21a4rkwtbYBxp/QglZRQGjjsQicGb4ABn7T6qD1RXgf3xIGe2yjQ2nZaZ
daL2TU2LET6lT4HpLgTcht4/jbvms8dHy5MOMnSgSMlWGeUOm9aR1dfWUYaHdB5Siki4S04xNCjd
p0ijRMoGsS8VlFj1FFxfuSDo2rR8CPs0t/szqPYHFA/MEFvpdxfsAIGaIZ1u/O6qitSgHM+s6JL3
41kB84Y+he+P0YWLpEl0pNZkRRIu9jbfSfq5xxxScQghId7MBJf8yg8f9Q9duFJUEn54VXE11F+7
ChWRoYWBwwot7oqAzpR3omPr3MAU+I56XqBA6VziYmfdqI/cQGRlkhMk2QTAaJPepdEmCblRYYXs
xwMFAypz7jCvFcri6sKYf/wRRNXpJMyCFv51f/WNCgoDh4LK+qkW5yrpCjILKFvx1z5PRvxoRX0T
5jiRAaL77dUBRhMeaRul1Cdp00w2Qd2+8CBJySdO+p2hHfvDnp3C9hgH0+9HWnhipgzAJwgj4YbI
7/GtueY9HUHzX+mcFp/pc8A6vqQkomp9/CfYTmcUTX+KtDEqmIY0wOfhbDJwI0ijNOdYM89fTag4
WU9J4xzilvdxqLCNWL8Owot2DL6eGV5jK3kYadtfHxeHN+abRBjJMIYtKI/mZ7q7+VC91xJ1XIjg
/M/HoifQU1zo1Hc+JRQ1XWrbfEbVu1xNtCZL5JU3XTDgVsVvRsANVjTrDCToXvoxmQP0TbxllCxR
3wqYx0nGERQYpPliZtZ6lBnVRqdHxEgDGOrfyC16xlX+kZrlJfhjGzTDe8CDGqFR8ZHR9AQJeyaI
gvMS4QnckzdoKgoAq/zC//WjCiTVWwMYRfR3N7iQXtPJgRm26h7dhpDb6sURhI9FljsM+ZuMeur1
oAgdnY8RWUjPnShjmoeWfE+0uET1oJXX4NKtv2yxb4icHozQHfdjx1kWEVD4DItRndiuE4ZgXght
XrzrsBcetXi7MBFnUL2hCEpjDX3QIq/xf/A2m7tuAN/mcr25iCuYr7hUM94SiOYiPd+j7RpXo0Ax
lv3bXzo840B+sBZxZJrvekLhVLgLkeAPKc2bJPhT3M5WYWXAn27S2+PppYHKHmVUuw7MkwSig7g5
yGcgIrgrGK2RK/PQmgHSiV+fRTIHeCen3NjtdtX5ElvaJeD9rav5VHETk1u83LcPJFHMStTkN8ET
h0nNelB4EP+e0IdnMIn8GEfU/tPi2fA9W1jO5FpnXbaJ0SCnTcQS7Uscl23i0Fw1oqe25KIKFoSV
m8TKO2bSo8ZC6ddRhZ4TEMCrZqqIjtvuc0tk8iXqPKad943s9YDydpo00fju3B7FH93HqTR3+znh
8y8uCHr02q+i/bmSjgTrdiU+2kyJXn+Xf+HkQSokPt75BcEO5YMwhvpnVL2VlJWGZfdnjFRZm5DZ
7KX7RSzyiXB8Py0xzFbqOHweWVBu9lL68KZ+aYxSMr8XIsSzpLnJf+3ZsolD6NYLzcv02nLBamQB
7pELq/QblJw0aJenXjHSSxnnyDEtPVelRwkV6aeFH/9VAX6v3wDtKXWNA0S16Cq5fMPGSug5DjC+
qsBufFW4NtXDn+KyIlRrbvrq3V/Xsd1pXbGgoXrEmDGLJAdlkX2GoNsvfoldBVgJvV+r++CnTvSr
IQ3xPLY9UAQtETQwHTdcFnVnSqBrEQmKKWRFNQzFFMGpwMCG5qc3R1V4n8DPoBiU2k3+8nXmiAGp
3Jlk7MnW/T0gX9WtccrwjSzXWBywDbchn6opB1PY9ebyFK1/auh7yiFRGFqqwXdRLtTuGW6s9p7r
lOoBlUborOOtTHLp3LaBbkr6qIBi1pQ7uFdrEID0hVkh9PPp9324r+7LmeO0I8fy9uKDWWna3UD7
KIj30wFkeCz+8Oc4POExbbdzS7I+aFFntngIT2M4tqj5cMQqhnK8nVViIfX9qEWCHaY6iCPBflIR
hxgbF33LFLk86Tdc+YFe9Nguw2TxGrVlZwSlEq9jE26mtq6Qkft8xsFgINKRPKCtg7bcUu/zaydY
k2PzeD8Hj5MOEL3vMCcJ36WKP4hwX2ue+IdECZQMW697SFmfJnVS25Fn9h+aWwA+I/lYM6mjeX7i
EfKuG3kGlpOlGwuhR5U88T3SUyGcpRvO8ggJVe6jJ4d7LjA7CVvntCbm7pbms1CB1ujritjy4wCt
3G1KUFaAE2XtdICtNvKFhvyZXxIKkYxo7GZcFyRkB+hD2Pyb+SUcmT/HMZwkiUBkyoSqaiO+KXu0
aPPMIEkeXHeVNEygvnqnRg4LMSxiYTjfRiqo+1DK+4QI3ipKss8hzgcS9/gdmEY64CrfLlxg/q82
fKp9WAETBI0YOe5msaBMlvsxMnLQWct4RVfyMP10pUk2LjgNin3JxijjO2jkrEIxQ1SGa/XvV6st
3CAbiMgWrJqw2/DAWvD9w+Lk2QDYr4EGcEBaNLpw0twzQ8E0N4BMLx9T14BQmr1znsXI2CS8rwYM
EaKBv1+dFncmeEDWI49BrYjPxeCGg03TS3PLvz4Tr9oL75ZkaVPMoMYpqq0fu8hKrtKU7nFavVTN
6o6KNkgoag6F6zJgSUW56qAJr2nfi5jnDdizYqFvE6vhQsH/6zj47h4r+o4uz9mo4jY5WYDPW8lj
DzAa8g7FPVnMv3qLasWfGGDb7UsPDkMXxwTpaS1YQ0HStDO3Dh8Uz0ozT9F3Hq8UqhXqNbi+7jQk
SB8kiHuowEpXah1V7nzPgl4FyerXd2yogQeCbNCzLA0+aUdrGY/AJAQ+9Ybpbk3YiEKdwmh9iI+6
z7oUWZK8OP4RL49x0J8ysejaBNKsZKDD/6TEJC31OlbcIzUniawYpMTAFPMpQYhmN3PifGZkhGC9
jywy4Mjaq2BXfMNQU4XRLVwmySJDTjgZvwZRqJl7tMyH7r0cK3Nj6YJ1tTLbiLylJOwAa4OI0GMP
DmIg/pDOjFL87IAR1JnFtFmqUlodwrBCuRzwZXQoQRk4JfUwUngxzGiAhxw27E7s1FNpfyJWJlR6
0A9H7kyS+jXiS4IU6mFXexYVBNUykovCUDIQ5ZpujFGA5ACw5Z2ehNJyjPpqVM9yUhYcnGQpP0wB
lURduvpsm5pei4eb7wvIV4wddTwyEC2x/Th7IfoA6FOwbvySDwJ7MXGR0Y3t3/Lzsaogxu2Ywel3
oPA1hZ5bJps09blas/EnB4/N/Z9SZprAONnMql5bARvT6TDNbf9QUfrp1v/C3XWLTOINzeaLvKB5
DRa7n0zwSWEngoVVtIAOX3EODtXHw3O3gVZXloyV8eTvEn5c9vzvLp3chHmxZL0EdY/W5hxAFAwx
QOJQT6CAn1AmK5DNezJ9Xes6nvZROnbQK0igaZRFlJuvcTwn1DDbpOF8UlH2omLg92CBPAqPyPo4
BP1XFbBT0TWBPDmwb5VMbnuAGhcaaJ4Y1iMWXZxykKI8mD+uPrVcnsqeM4OkKGLTrr170UbDV6i/
xLo/5ovUx7+++tpbKYHtAE5/K1gkFCBuHzM5vGPcBiNslFsz3TDS8wXZBRI715MgaOggknfNqJ8P
4TrNj/nQBy/cXhrB8bisXlGO1ao5H7pQF71QUF4AFvh5eKkGIeK0CrknJO8VLunr3SBEzGd/uERR
PlMYEnQnMs095sG27Q91kPYK8kY9tKuBpVkGQ3koEQ0ohgUtoSlNoslkrzlqbPIP9UipwWg0Q3GY
1TtA26oNrkOOmy0+CS27o0LCjEDYLu/vWYnMtcvSRCkt9H4NAz3oyheU67YNczLldpgs2Rr0u6A2
q4ZpgwTJzd9wm/9gr9aA0EyQ7+cv/z2aajmhdF6L0aEg/gTg09OtGcBkmq11tOvpdEzYdnVBrmQQ
JiU2BdCWMKVvG0s8uZqtXZU5X/775OIG3u5xnzNfYXLO6iupCH5gzWWUcPkaf3UNeUxY+irvAsxi
oYcaUKywrjXgYUb4pZ/SF7ySSX5uRYulJIhJ+kUqPkbLOR+TI0QLf2YQzrtkRVTIxRnb283mkpIe
fVaO+msRSfk03/bPwekcsuUpZhDnQ1xBKRXa98FNaQCSrGpT0xGVyWz+LUZgjQlqP9C7VAkciVuX
Rt2MpKxbbkJi8hXoFDLDNPfeaEJB0BZvAm0holXAUAk+GSxZF1d4RyDKYhTRBQfWaiOwS4pNXJ9e
/JvGxeMuXwObUpA4AS6YrVuJ0xrTnrI2SNGTNMRU4fbgVhoQ5R77MinwcGLnI/zIwh7SQTr0fyiY
QJtHjbpsE1fUufDWCvktUubbjrOgFt+ZZH8gbntkaVPG+B6Q2xTOKG7R490r7R4I3xaMmFuiRdOY
Q0Y0eqJ3ncuTiH1LaZIIkkwoy0lxaymxiYXOrKtqiDQSS33fRNeyS8uVSrInI4Bp74lNTwUtOSIA
wiSoWszRNmO2atukaPjMLs8K2pas5I+DRHkcKEw5FatEjxk1ElV9krRhXXCw8d1zWwjW2L/a1FC0
GJHpsobWhxaYroyP1MQnmTNHb1evaEf98A2iamK0CwyUL1A+LVPIHLxbx5egRoPtJshLxZQ9IfY0
5VbN6KZJmEdPPHAIhxsQWSNn52J1M2Y37wFYSX1uE7X/HEOifQQGagVlhVLuf/Gyxxs+TndsJrNe
5eZrDWOGpzk3MFb1e/rbATK3xhEdR2HYR+4T3iU59RyCpn32Shu8w0kg7t9RHj17S9DYHLyBtrTQ
i9Qv4Vo5gfNkcA7+fFGMhLXV5tFIXOcHpW3fe+diejfYgmuiWeSWqa4AKP1kVySdsmkUMN716NLP
ZYA17sewURJ/o/EI2KKGMNuDaLvcuQmMmpzaZhz+0Te+Kdw8Lq6jKi+JcNd3cLhj7TdUTBfcz+Le
ZbWdQBXutJcwXM7xGyuXTyrEbGnj9TLWFHZFFbk9q9qszxQQnMz4J8yR33/sMRnl9H+JJkC3R69e
Amnc73C+NTOau/1uup6bcrgV9wYwnibA1JhLua7z6VoLDSxJmlikd7X5DP7CB/U3YVHvwcX1I+7N
ZVU7dYgNYMmKihpc2tN4YQFvSpxOKVOB2kiU2ZQpyFaggTlzH8OEUs1jKoxxDR5UnODwX1DiG/DS
nGlpSVljt5DgebqPAP3+/aubHcyEQtwFp1y87R5I0RHXMAhHTEIVMxsuqXbB9ag7yb880JJDKBbe
HsdEBQ6m+TNSoQ38sOMGqYqlNGBGbFZNik6OLOiWPWKRnl3jRhwNHrYwfL/QbhDuVcWjWQyjzRJM
CRCcs3vBOpmPMOFhjRMzrmiCG3y9Tn6k+1BL6E6xh6eWsWYe7BxoMD4JZ1aya6GcXYfIfhXfPDPu
+PWajepiOsLX7OEDwJZdiLDz1yayYx36y8XCrnmq+xV6TgGdvTAyTSMREURFSCKU6XGQ8DY0N4PL
2CFvEvrPnPU0e/T4suhN+/MfKRIKJGM6rCSloQaIeK/81E639YUWnY7fBbCi3tXlKu27TC43jqOg
5bYe94P0R9011BhV21qa8Ftd4wsX+T2xazQ9DemOadJTKeIaq52kYkWtbWiEeFwLvPnsF4Hko05r
FsmFmEe5+3ByaYBJAQjAwEaVhQBSpBlX2Oe2ef4HC0bzNYtZhN8glAbCirOnzsjDuUsDHiKjWu/S
o84tUNONCOma5G4B+FqqWyxWulRWdPM+h+xfp5tV6WHvDUTw6pcviYoemuTxmQnLQtQYD7fs5nqp
S3UueCPm37eWwHiytrV1corpzdbC5ViWyMOXn5+TUrMaGaqWhSrUoGqPZQq2SYOE5m6gCYQPtOBV
GnXfQJG8puDzlTHv25L6fvch0Py3MoScLat8O8t67aFYo8o06E0FfDS4eRchBMRG75vPNAyltumx
8GyK6WSBZC6Y89CszXHqDeUNqfKDvLoG8kAK7ri1pqnyWSbVYrqa5hfV+y1v+naE6vkl7ZbhcJ43
Jt3RptrsJryaLz3e/8Q5sYF5t0MxPor3a78FM0Lmk/i7+9bn9XxfQCrzMD/Dgpj0KuZbRpX7WnRD
gvh8e0eo1I5MauX+kl2Z4TldMCbx5AvzVGFuaDt0mSsLtHZSodkRiQDUK6F9OhITkePxgvbRhI5H
Olo2XTvrEkcxIHNEDtsFHM4GMQzHT09BbgYL+6RRS78t9V7/OU9tJlhNo2ELF/AddXaNrISaYTiH
92TUuU8eTSSFgacqQWYvtDEYnCcvclhriyX2w+dmPWpb0pLyw1tNPYbbxaTDSRwivMaXX1TxtYjg
e5ves+rIge9YxBXBx9Ub0RNm77l1MpsSpcyk0BFTqx+9UQy6si+she6Va/6d+9HgOuYMRl+kimo9
cb519oD9weQ/UYjtM0JQQKUh8RQBzntKoZx29nxVNbqYxpxf83TS3nm+M8Mmp5Smjk9EgHv09ydy
egKiS+m/tr+Ja3yQukfaEWDW5RSuiS4RzmIDJIvpDemRihLhxVUevRgbIwbVz57+aU5MmwZXzUzB
g+fjnl3QSUCjmlIJe65rZdmLQmqSVKl5L3rmskC8Xm2lEqrKAzKBAFkmOdGwOSE6pZGKvwZ0ke6x
+DkQoNUpYhncFWsM05q2TVtqBNmMFeb9+Huvow2eNUkQG4TrqTyu7YvANv/ezErTPlWg8O4G5tRu
gV5u9/IX9hydKnL1B8SWNsp8tZY4a6gUMgJr2gLvhaOpBtdp0mNrbWzkfIfWl5chExTcm4EwDM5e
TcMAoZ7Lhd23PnTz6RNs2wC67lMb1ovnVLwm/FveC7JoOmMvT8YqN+v3YEeMpXNfk3Tom7OOYUgy
trUgn+QEyl14egLqyF3Tyafp5AKCqzy/ZVFzmDCo2mSeYg/Hx0KK2UrhO4mqsF1/1IH+Nm9vEObh
Ty7nYmDZJyUOFc01WABXVknHLqLMu+ThswYnh3SMdiHu/1/uypdPVsqCxTPOw4RkLAZMXMvMY9Jc
bIm/1IL58f5Gw18yZe6CWjNqCVBLXBoz5dGxX6uRp+Atr50tPlXIZ+1kt/jKUu+C9aNNmzc2+56C
+H2odUfGc2Hdr6BdYc6yGAqFOKH3LPK33KOsF80c9oSECmTWYg0dcNDTRH9I9+ywypT4ShJ8QMP5
WqC0zA4zBBTxRFD/t4ST6nZjgQ+/poj6hTuxLqdhgIOBs6TurCW1V8f8uSaPDMowDdlabjBlnIrL
Vy9U0cSV1QMo1gSjxcrZAgbxYZTqfNMWxkZIKu1IO+Ci2ekCESkJT/PTnwd3NIQyb7fx7UuroCkK
oRzb99mlIskcjugwYMpvaQpvNCYUrptAUWUITxGI1FatZt4mw3lFxRI/yolZMNdxHxaMmwiZ16ca
rxbMm9n0T9ntKf7Blh/58YdPbpBSXhFe9ScP7nNIY75jGqlKLKCbnrGvtskUHGSzq3rsjwUO62gb
ccgmLRceOLCLGawp4sK6BMTPchhWt/O6/w47NKcg52qD+LHBeQ7aRoN28cfsgL0lDAqRIO4XZMwM
VxMgG8n41nr2ObuvSSon9jjZUVk9ZezqARV/JH8yJnb/qPDC+BVOVlNzDXK3RtqjrvDz8CAloD5O
pdHjFx1+95nyYblXUpmHXY7JJQdGB0vYIHj9cM+MF0I3zyhlZwf2VBVdZSQLCOzzGNJd2LSbk9xu
8/Ox9zv3nSp5rtLR3ZLdMypIjmQDhR/Hqx2HN+aJIZXjbC+mKhWvV0xo61BFyxFxOzb+KgOz1F+k
0l7o3qq9aWgj5SVn2L/8gFdWSsRuVSEDoAlJP9JCxS1rHa4biHo2lRbLlfR1xesUb0xmlyU0B5M0
/I4qGy0h1U4Fqvou62s79J2pQ/C0jBx7S3bt1V+GMTLipfb/fClUwGep5exDiYkrQRNUXDdGpatK
CI3KU0J9jbrX5Lu9v8K4kvp1pQP5NXpDVePxLIxLVfIGjGpFI2PPNmCADrZPE4+7xYiYDSOOHmuq
MT0055vM5jTJ7DbnjxNU2wolOV1dksmSMobfL2UdWEncizupnB9tmC6Tlx5E9XpYVkFdNbeHpQ3x
hqiFaJLWnQLuwNBxeBEXWITNZd7wV/XHrL68L/4o63sa29kqfNf6ykJ9M4miNcdtR7L1Caw4Rgjw
1tBemlwGI5o66YxW3zQfhAg28n7JTePSjwiJ2ycKu6EuFevghxRWSk9Lkqo1/1zcsXmdIw8vkFln
tInuVmUfIDObZ53xnxjN/yXVtN38GrYZ4+45K/0O41RA9PL7WYJRFJhcz2Z9SkGJs1c0peYJq6zC
yGoCw68zCk4XMHULR4oZh7GJ16IkBcyO1W6cq/7WWWSZGYXKn4gNbClc5w6B+e8k/029pBPuJezl
BoRbWA5mZKwd/b7GD0wQQwkTXYFvlPMJgwKN7lIO+Z/gqMGnxu0ynib1h6ApEXrRsKjQOWw73f94
XL66taSMUFsYKhuFiP09qi5bqyRXE7YHIT/AYkv+uaz0jVLM81Xjp92WviV2FfVLApWcusClwia1
F6R7RqbW3bdn31frm22RhvsKSVXyOpVYKfwqwRtarhfN0h8hMTYhb3Z6hPr4m92EffhSV3f93GGj
L2W1R0KOYmInTGvN8Nxeu8ERjxXtiR42fPzYk7/+wQq1L7rDNbr4zBvNVVYAG2Yu3A/PaRp0AMAc
g0VPXFJ4NvslljB1OjVP1orp3e4uewMnUrmRm3IF2sD8dmYsbr27A8gSx78UNEIExxnXTppt9yMq
WT596BuySgyVhkTFh4vxDmGca4ARvHduEHVvA63OZSw7ZG9T2tTTcHQpMrarzVmLYN05h9G1xVzy
wqqsTXhSuYbt6kiroowk0OnWSkEZclIoxs2yQ6XTinNeDiXm9eP2CW6vFpBygqMT10iJ+rSrY/F3
h7kF8gDpJ8QsSvhHlfAC/m773HSe7BEcnYqGvzJcnHka1+oFXXqxBOWYXC3O0intJz+4HLz3plja
mVcrnOiwZpLLKfZvhOOcNEvEfMG+GAd9Bdny8HvY2GgGST+WfMZteakowHrpfAsZd1QxcnGD+6Aw
TIh+NKBUFosFiMkTW4O8kQey3ChzcQ4cAJRORHnMHae9i730SZlb5BzqdBcS9p3aXAQXdehQSwMM
7sNMzlhoJ2eLW4PcAJQMjZeABP6ZoYcsd/LVrmDBNQjYWnQaoYzSL9whQdXne+WXJsmY8LppKK2D
LHPHKrpCBcaHd7K41PFNigozLkV1Ks2RyeTs36EMz1zHMJWo/y14T9DnTHBmHajT3APabWYGuV8s
p5xrChxnE4ew7DmUg4DPztrs0LRv0/GAVqkmxqxe/a+mwL1rqD5B31Lh56X/RKtvc+KokTypOvPj
eca26UYYEGm5k11TDJYOV+TjkcXgIEG/P0tzKkIV1vmxbRBGnzW4udmMylLz2+nxjMS9ezEknxzU
7euwg4Q03oM4PL20mGupPl9giLBcGAB5lE+kqu8uIS10zE5RSDEtIM0R2LKj7jTOj1bnHVs85dZd
XJkeUQenRakxWz7zwVNYeA5S4XijVAdbMxe5f0nKtf4X9YZRDtgBGpF8XWVbDmnU5SDH9qrUAZl0
GOO8L52XmfLlEOU76JbUWzeuQEKzr/gbMi9wttxnPaCdnAH3aIByQssfVTddlJxLgF1puOyFB4PR
AHm0xsv6QrqKbLe+yIjjozNkpemYy0lWp/ZV5NHz9Qnd3Bj7OAQ2mUxaizlPsTP0MHUO98POOul2
WD6eAkoo11cItiliXxBHdIcdZR/XqpWusxSvl+rtZpzvimR8pkrAYRQSfqlZZMVuFgDrH9tWfqko
ro64dG4SFn13MWz4fBPqdOAybEofagPsZA5oSHGciQBfpnU9Z2TdiBFnaAI/6so9B+jWKMP4yI+I
GVhXHXkySxjIMGCMvqcfz9zyQ0QHoTn3RtEtDolj2FnWS36sLqcafH9181onqi4VqmSwFK92uP2h
4VP/uO+/i77ceQTSVctwJGc3SXGda+2IVVEVMop/P2b7Whm8FfHehxkhDMbqCZLVnEuEuvlgoXi4
ooDRK2teHWIeOmj5mq7zKoYB6CYWH8U/PnbC2svB6LRt7IslrNjiU2SsuI4QsFXvxE4lAVPjezaG
ojwhH/Rt1ruyPP1DmOZFnajjIRtip4FFGkhDEd6Q9+Sv73ihZatN+fPdvaF8aA30KFTnPapGDI5/
9SGMWWBqZfW4tnrTdplbAlgXee3/t11P8lZ35uKy5hn4oQO8R7x+/Vkpv0CDh43awK3JlESBkJV0
fPgLkGwnjT3X986yMQj/FdPpvmwbBht3hQGurAlNNwq2sGTuu5FerQmvzcmC0N7qB+m3MKrVTN8w
/otn/io/vslrPZS6P3if/Wl/K2IApHYfNYScoIHchYjNTyE+USmdzyJo7JJzAW7nHu4WKt//PDsy
aXLEhCOj9e/ecz2F82RnEYJAOke11TYEQhMOwhgBpZ1Dk+MOHEkz+srp+eSRPuhO1DK6n0iig88l
ewP0ngtZ/oj68taTpCRLsPMlGbyaWicMpyP9RN+QGrllbRWJusb/TZfLIFUtOVeQoonbnYaZpOCN
6AGzC5eq+XX5U6CYbg0OKj6TiUCqqOUcK7BKDufBw723HE8YuEtiTuozK+jzfUS7kqbDRNdkdUUr
Tl7bPhQ3qxwUvAVN3KXrU7fDiX+EcSAAQKi5964vPuTqDc1v4wVLYPikTsynnEhOW8m1/cMruY4s
TpY5t64F8+UbXF/DXWcCxFP6RyqATpal23u/udqbuDkWmvRtqug4oxkKNK1HLHHV6ocPci4F8T/q
NPbamQs7jBWPIy84Lwi9Qg/Sszoi/yy2cDkdIgw80b2BGwc2IsZV4iUQQh2L6y5EuayUH3cx33lV
QajF1SH7IRkwCvl+BLUkRt4qq4QtZidFqFsDiK0x1Tb23js5Nb7nLcTErvKMPLH+Xdcf4g9McHT5
/heEXXEXvLhmqSCJNbc3Z95MC6jQUYshMTSP+cgsXjjUYv4CbHloXtnizd0UcGtqjsg/5LSKRoJb
lMvAeydO3hz3iWIwh1qF5nlhC2P4dOjY5J2Guuiq6718lPe0MQGzfr28yb6FP2GzAX8mNXFhRTx/
X3sYjkNMUHneIRtVsS+KEUkE+Wca1NKelKbGKzwaFyall+AG0WKT+NZ6sExlMWzDewYbxDRa6wQl
xzqHBCbsLok5+irUKIaeI5gzsuk7dixMNeUqtOqIfp7LTtJmjkyhtSpaO9q3v/TsHosLqlvJDvpG
SnUU9qHDcQU215HT/Gf+Zw7iuqNHXqT0TRnYfK/VAhZTJetIpW6tz5w95mfPkGXOAkL1XB3/un7D
AxRGH7Foj6KXK8MUJC0j9xhsJqTBG5D87hEVo/78sR9OlNLUraElA67DAWNHK5nWyTuC1a77GBX5
EFug4NT1nHD5eU8g2HVxJjjmwXmuvkA9LQFGYFJmkfM5Lvs7QCTCxLhS8zXJZ/XQJEWJSnYT1dwo
m33h9BYWTWMG1pxrMtP9NFgskpQTX+++e71ef5gf9qcj/y0n2yPf+X86sYQw8xR/zjkB8DFK9WXz
/RXGDvMobB6f21p1M1RBXHMaa0Pz2Pm4NoxzQcP6Try/FUbTsSyJGj1diw1takbDkgvv3Q/p4+lb
jMKF8E48KCjYNTbSvFpIaImdHTn5CcWVyHsxy8eaWX/ewgSa0WgHOoopkoHRBrFRSLimEtinKKBP
8hdMJvyOuskKBfP872M8be7xwvRbHrvJ/qMvdaJ7Fr9Qv1QT8I+XIn4Q8iem1C56ckj59CM9ujkR
S4i3Bkb9s0yBjM6cXjjL+fEipfmgJTy1EH+afSYY+UCM6fjna/0h2DVNRty5W2h8+Z44i9U1EHqt
tN0V+jELyAd1UzUW96LjaqtwXlqKo0lR9WKOcBbabht5SYxqs4ACSmXGyURClVGtckXtqje+nPS3
2daeHNeU4JBCwqXMrEqnoyBK+fIAUJi3+u9Qq+XScgE20+gbd1ADqHyjaQl1QVusv0Xlu/h2oDjQ
4PaHA3wpxf/mNLSuzjDwc/3djdZTtPs8fQAHJnYYTlXrImOktjkuMiNTlLjwZI8azzII7IfkHghx
JYssF8J2bMkmvOmKr364CKELdBKWnXiatylSqwcPwGQwigQEnoJaYZdDUR8qT4ev7X853ly/4Cyx
Btjw9DBTxBex27qDFwutjLTQ+mvS8VKTIObvH2BAjcyLJWZtUKNjDPiVzKQXJhSpPcKD6QOb/iaM
S82e8aqv5yAfm0i0iC+M7IraYfSvDkFGDSKpxYrAivm1A6WPb47W52bLUYU5ic7n7EnBQOdfRZih
1OCKoY84WTg96eNZ6k6XEUx0wXRL2Sb25E8qVmOH+JI11LCOpYo8mCjGhAGRyJTqVQ/jwBpKuNSE
lLAP/Li9u5QzHFNrOdAR15eM6bRmYg4WJ4pG54/AaTqvnP2nAAHjuZ/a9IJEoVmuHdKad8ZlU5lR
5DSyvDTggP0m21wGnxh9sTsJpJPu+Pn0mlLujfL8Aeq8okbARASEycUE3b6iv5dwpekZI5ogWnDW
1nVnEEV70UcfZqfQWQOaPqEercf9UYMEYChs/0AUx8Hf3ZoMbVUrWGJGtC2tT3KTK9yAr2YMG3kx
3hU6NcT7QVDKc9+M5Mln05VBXY1zcvv4qvw0m5Xb15NeCjKK5FtKX/+vvI5j4PzL72FCkmtz55gW
4UuYWX5fKnsOybozf2mmJnijEjHQKmyfcJBEWB4s+96IB1NRb8ohO7R0OufnYw5NLrK1leSivk1H
pM0OFF/yfdL8CU7NNFENJIa+TRZRj4he627nJgXx/MMsnXp3GV69yB+IajH/v4B1lwN0/hrUaZKd
DVFJEKS/TzmXnYkjGbzlchVpTg48BduUuGGWWox2M45sMpWx8dV7qjgY91di+AhZP3TO8rS5dTgT
mdl+YYwXRtPRqkIdjrMPDhymV9tyle6pcapBA/OSD4x8q9PFZuL0hm4CMzXynkRkY87NnEygnubC
CkE4Q0MRgKq9PTXKJz8MUPSNp9wwaC/rSucDR5foFNUfnl/RexGP52r5MEncHjmt7J7tkwKaqBU9
gtzzUjZ2p2ZUzMkuAQWxeqd2zPvntXD32il3VGrftaN0PQyz+IHmrXBUHbaVhDKBT2dWeXoXncmA
cbcKx/6CHgGWfDEOPiWOendLrsHwYZ2bA1gf1kXNBKvZwvzKtJdxMxhZmXo5b0UuOMDnsqeAMlcv
fXrEPzOiR3g8hfPd8OZ9oZPANPzoyQtMZq6lTb5H3/4j6tin9ltb4N+M04FmunUGCxZYAYpJhzmb
fnAjN5C5VLjCj7qfyl2kGvgSgwl/bH0osPEoEL2fFGP8X05c/SzfHsKEAmdXoPkPqh1Zn4Z8vMio
HLYGOiMl43Xm2PQZoTT1h3KBpR2VYqTs/GjcA0l3xT2RDLk7eDRTGIGuQNfueE8F5QIfkP86HUbE
01UcO6UTMsH2tpTvR4/RMvAr1cAxHH1qrVLpkAzs7qUDjaK3i2djIcB6pHu6yIQ567SiMCP9MHmw
DpP5EtF5RDMpJvFD6wEEwkYwNyOwV/p43bwXH1Q2zolxUFJkJCJB9/3vVD0jv1s4jUUmGrXeYYqR
c/jumdxlVPLG60246zNrqL/rmlXxzJjlHKVRAy/aG3ZBiQQ0AIbpl1UDxK7usiYsTZSDXlRxzFkB
RGeqg8uiMDp7XJvfdUu3JjKAcsHXY03oDtULHj/1/yfM8xhyX3wiWLg++O6mHPcQNprSiBL8H58u
r7vdOKXm7Issyqh79bZT6AUZe76h6/B6M4CuW1bEJIN20bIYgtuCZOQ6Arx95E/eyf355oOFxiG7
vsBZw+i2rrVRIvijs5a6kdFwSqOTPR+TgCXe1Jy0Zt3p/aTzxBYFdItJAWsnvrnHz3bb0/jXJLGb
BqCtSJrT1KpB0KCpWGCFw4YNoz/uLz8QT0edOQaoGFCKP/cF09oQD2SvuV6PyzvFOFOUxZS8LhC+
0RLaNPSCn0lVII3MV4C9rhjnQSYeV10/uPfeLmzy7TPOsMtONUBX4iytDgPQE36Iw3QmyXb/jPlt
Qetu2adhi6vT4P7sLreUf6V4DqpUQKVv2yxpXqS/VCrq2tnxhgYQy9PZb2+5hnkDtLOWX5bMtbmh
yC8K0fwm1tt2xOKnSfsOE+OgDhSkbC7l7rnCR3FQdvMmk/XDRy4jalTWQgcRJZMw6dhGMN8KRFDZ
vgJJlLMzXXwkWWc1eRGTxg1Gjji2XgeFuxqc4MtWc0hHzvGgkY0coeYRiMgjgRfvC958KH53NntV
dYZ4JllNFr3YqVnZ+p0C4nuBqqD9RBgzaEkM1VXXg+id/nERHIvHfMm7onIuSJPeEtrEz9cDe0jA
aRXSL+GNSpmvqGqXFTKQF2EFJzwOvR5u7bTK2ybBikTj1ePWDJ7VmOelK3fPSvJ+l08kcNwnrv0U
u7SD3/fJOMxxMD6HxXDSMFwoIx0YuqfrMDdFFvGxmo5nw409QqylJZ9bA6fnxugs/Gb8IWcbGidk
PgUmFxbgoM3KXrzFhI7v8N2cNG4WAEDMcN0hfFQ6SBls/IdY891VTOJbsxvu14u/PD8B31FMFC8I
Nt5VSb7WBxyGQpJ/bN/JWLRAsQ05pyI8vP8Ooli+Va4+m7rhZ/CignOZ/F6nOuehHVJGWrw5GBl8
L20V+hORQcec0rW0uvFEbgYQ2ehIrWdFWPcZtqJ9eImuw1pVNBD8vUYPioJ6Jw905U9gzTTt0i/S
MHe6oSSjBw5mVYTwAyHSYkWFh4mlOWh5A949XUCptRsVJ+dTfyIGsL90WrZnL8xnxsEIy2jnHnkq
yGTQB0jk8Tkil8Mkeb/hEx31I9kuAS8LOeFg/Ae/OBivmxNlV+6SCzgTO8xNIKC8MfYrAdHQU2Rz
ykn2Hp5PSPP+D5hlh4GywiufE02oRuf3st0gy5o6F6w0DEM/OQLNzQpw5lMMwJbVWFAixWxBiIXf
821ockW/wXycqIkNH+P3SXH+QR/vo9e78nNrIKANrG7ud6qAPbVScZO+zQ77ZYifjm1CFUCH+VTL
jvgO1PkFetGKtOB94Yp8cUM18b2N6rpvQhC1IOqG9ovoWP5P91RMwcI81aw8zGojA5JlVitYuyQc
cgpXhJNG6yt5kLUVEORWyxzXrxeXsXJ5oqZNa07WEZCrYCqKvshFxRMGlsXF1bjZ1Eiqocc4BXrj
NtlNsZwKHbHT57nGzT2RmV29eEMca0yhcxYbPMrWf28ExgyVsog5SPjnKDpAMrZCyhZZvrKWwyLP
Sqv/GQN8RFmNr2J/tdnmsAfUmUifhrpLTh5U1QrBeN7mJccGxGtGq5yobeuynq5ri8oS80Q1oiSn
mDdae8wDJeNaOlshJsXOlkpDMbYD+hFrRHLp9BeBBS23ds6ewHHjqw/ZC195jTGKjhkv8S4dMa0+
mh2hI5lpEzKPTEBqMLxXz9ewtq25NJnpkCE0yTgssTEuYA0Jk2uODFtSCpLpRgoJ8EHJ54l7BuQS
wxI4hQCZOpNhGBsyUWZNeaXwaK5FxXSI2kphVkAojXTf1HG/q+LoRS6xSXY86v/F9WS6wkyvi7tl
UCfg9zR5ZsgVIAuo3/V7IB2sm84eLt/rqtplT56lM85UiNHML2mq4hxk4xwPSeWm4fRxyAYX+N+2
jlG47wrP3khTg2zRiJvd8jQf9bwohCnjOTb2SzdJ1X2UUlIW5LkWEZcSkjzE5cOvNxGLUX5nRfd+
XdKeqiXbb2fg6JF+XYHnOWmDf7YM/M7tD0YVp3VUELYMeUpQSm0aqqK81nbYUmFAAeuTl8q5hdfz
/LGln+T2b+TczgxBZdY5ZQMLxcyJBfD0oF5iLrfeY+PaMh3KvX5pf9t9aYroZllV1l/dYIPd5hHB
h2pf78YQyhg/MBY0n2joq4FLXvx4gXU9yk/k2/J7Jgv4UAmpneMCIjexat31GUL2KwXUX6WBYdMp
7NxjIrNojrpOP0XEuC0Jdhs/cLBKV4NB5HN5NM6P7GYutUBTk8PYy/4r+YqQfOVauCfFU8gTKYKJ
SmwXyCJKULY/UmuqPkUBMa4WhRM0QZCVXroW6fJXifwA3Sa1bFZtJSsojQdVBUBo0gG6SIok2u1v
zUyKatPDWjMJVqNAGbQ45+o7qiTqurAEitfrc/E2ZVRFwxH0OjAqv9EBYM54S2AAmHSFV92a1BLH
U32ORATGoPZXey1mO2YMfP56TMpAKh6AykLAVHbRQsb0WRcZY0eiYOjFyynG5zwAklvCTX/+OkiT
75X9YI5ac6VWXywNrghszrlHB1jS1IpyClwLUfmHdS7v+e9rWLFQdgi7A6qOYN2NWHuoubps5vJ0
cX9FDcGP7bDWGaM73MZmbliXJCf/IGv47miOXafYtGtoXXlfF+YzQo0h9v3/+uBJeenVA0jX0PbL
USX0rmPkezeCTT+1r6HxpDvE+/a5ZIiJeIfnFLY9wUgCJsMbP/Tct/eyH06ZOZiBRmeE53ernyGU
ncPZKlgPtAR5ZfLdV63YPv1f8CuX65JVOdesDu7c4YqNKYQStiuZXezP43P5rCEe4dmSmTwzbO3H
FNphTpPRik+ITlDU1DN27b7Zl+8dpAR4wr7MwkuG3bJglN4MwkY3Ebqq9daMsjG2HHCIMhXr2DpF
lzfjAkrbCWYc3+Iu3fsjvi+euRAZ6b51WLkz1DH2aDZJVhPugj4HWilxxVL/UxXJAb9LjhqQR5mq
/UaEMxug+8gs9lfM7NdBrAlb7KbBhCNBRO985MZ6X2oMgqBwSJ6+XZknfuAtgymCH/mkWFA3t68P
UK7ArJkjPbUKAs+DtcusPoA6oFWjoIQamvWqiyJxSuwPWOjHacUc8aL3KQOYt46xSDewj4D6qbBf
YRpZ1nihr9FXL0SzTCaZ0R/J0K5os+KP2QCjyMwypsbot8x4oaAqKTIPZKyN1uN8TZKiCpgICkzQ
a/sbpgAs2nsHpmDFguntzfUWn3obO2V+k8Rs8MOu7ADXccwsujyZuhXeW9m8HCgufahT4IlT854R
5P1taHuftYX6yp9+TwkpFAAfU7ABsF40tpdQvokxMxcK8/hRkA44cVSUnI6Wmn5etk/IOg3TX5h1
DexSqQ7d+YokjzPm/wcT0VyUylkUBeu7tXtxn10lxXrk1VXPcsAxTcrl5/GXudhPjtYQaLPXmw8J
jV6K4UDqfJVC7MRME5/eUbz9464y+QyjXoA+POmfQq/XHIFcECgGfHpANPlSBTQODXXF1bgh6ZuY
qiFnuh80q1v8WjavEwDooAIXS0WIa9UOc3g2/qaUnqIuJaA+zyGtf6fowqiw1fjKbjQZhm6RC5Rm
mO2BWVYgVecxs90nyKDvsqQevOhP9wMAfvjdG4sV5Op2lDDXfFteoCK76aWfVXJKqTSJiume2hyE
IZuodq9su/+7f9l8BbT5KesJGLqAMakPE75NXwQUgmDE7K/Z5Hvs9L3OyXoff4LdgMxoi0lzAMJw
xaDsksn4K1soNW9BjMvol4yph4H/Pes1mbifoe3cq3hdGTiUOXd5ZJRxlExgTs8rRM4UttmCbv0b
34DX1bE2uAajvM3t781H4E0ystE+EiqXp41VhJwzCSFHYGx4dqj7v5QGSHoWCVYkH49ps3hlMekl
DKjoJ8zFSrH1xkEQyqizmLc4z/rKP0+rBF9YS0au1qo2rfjUUjC+vx0bCY7qB3DtjJTvL3VDo1LO
BKBjEmsGls74zyC2xaeB93OHKloDssrd38Ev6unaWGZGTfuSj4b4krli0R+NaNS9omJY1bmxhQpi
slYZ/HaJeusZL5jUZtveopacoS+dkP/8Yh3wOr8q2OUcbmX2csVC9eTxe2GYnGVFB+PD/c+SEKi6
XN6w3AVYthKlmR3vbuoPtzWW5FKsWzshHvgDN9PhdjRORcjGjCp818HtEk2+nEzRd5kYxLgARtZI
qyYO5RQRpvh3xdGuf1D/LpCrup5GG5bSUm1Rmx1BkhHfjlzsyU2Y650mOSnJh1g93lO0h+OKf/OG
YVZlEJ5qXFAEteyX8vXXW2ufps0B7T0IVenvuKGv+uvi7SNOT9+hJm7lb40cXs+sTufHImQYb8rp
aB71WZ0dv4gbNCbzacH6gpzkpNEz9IKUp5JLeX/Uk92Q9dgK12mDQjRvfG5rAep9CMuJcXwAqjvC
b0UeHmPSJ0aAdaOzB4R78iYXKnux4uT2sk0zBQTT6geGfeQyMNOgMbq9sw4JkVEzPKFFvoj8Yk4d
WmVjoL5ob5e+7n7fXxcZ2x27pi2EZeerVjqec0pip/vPUwuimO38idyY/R33b5BkMsk35bZcNut9
aEj6VK1ADYkrwydwBq/y+pK0mMWiBr6LiPPw5hqULso1hkFFm6u939r38LAhvCFtITYPFPJuukgB
7Mlmi/j+xOz9n4eXFdxnEvdAwCujGh7UW82sujPxD83YkxNxfMQ0dm67VvFwXyHs5gndx2Rgg+AW
XsOYCFjbP2GCsHQrj94ody0cPFDF/TEKXA5BJAYAeQ3ZuKr6xttuZf2NVxo7EITQgQKH+FDdjWeR
B3oiBjAilgQTZATYsgIWo3/SMJwTVwpiikMIduFBr6j4U4YB0OIssvEjS2xr2RB4UTCa1wikGkP7
CO8CaYqxQz2jLnayqkKD3E8l7F0mcYKqXPVxCaGs4uq4pwle50mJ86aB2Jw6Wkz2r5LKiS4lIwBI
yySVaSgxXLVPLLzzsWmLfACwUIraA5YN9E6zFVUel+5xvmswqux1Uk0aQjGLk3MKDm+JZD29KbQ0
9GZsox0OhxeP4WCgLNpEkuecPaYpYLlZDkzHXlteVTlIVum4PRTbd+LC5xFdDMZB+xJrerO1Ojys
TQU3MD74+xAbcrcSImTkyzPN5r09XivQvPTGw6EBPhYpF31AZCUbo8extrVB8jGxPUQc0/3EAWGU
8/tAVRkJvM/FEulVvQaQUPveO+VLRg7HuitBITInb6Sd/omY+xIale2BuUzhaWh4N31HKHUB6ugQ
yF+nmLBwgAxOT2S80lNbu4d6SzVngBGhwQa22lWUupOD9JCBKwHEz+mavikWMc6pWBud90Y6Z7OI
/HEKeZ6cV1Eul49gBj++GZrFiyyEtelfqNZfTRgzndBCURHmx5z1PuLrwbD/dos/OQxkBbGxQ7kJ
VCKQgkATQ8CHKn5I7NeJOxDNKt72BCTH/+FGmty7PvBOVjuUm1TT88Vyy3SKR6jjjY4w6cXGQHpb
Rz+mZ2jsf0N6yWinswd2aB3mS5yZi3Epn489aLLCccnZ+6i0s1McbN4wVrNxVApu7DNCaRAdnq0c
E9X6AiDwLiOuwPiPHGHnvFOLyOGjzUFVtutiEiWATC4nbkMQHCWpy/Gwa0+RLmE1tIVPbJlqzFJr
QTzlW7hOA/sB/nzt9hbnk0zPPNKBYUDk8SPTSLTAyneb5soOEmKtLtjXHoK5XfpltxEQRho8oz4Z
/sEAxk2zxPyRgWxgr8ahjlGCmnMesDRX5lJ5ru9mTf7CBaIzozy+RyI4CPqiwsfYDS8XX2UNHkos
rmlE2hVXEusvcVxVR8cllgLUy+PqLOa2vXNYJjRjX4LhKnCA+N2AY00B2i82Pk2L78RdH2x4U2AG
s7JCBFFfLmTnVyQXDBHD/Fhv8J8J+5b1YxD2a0hPyXMWXrr7mzsH7QxsdZNAgPvvQkJprlEQObCV
lweIFJPoXLhm7xwX3sF87Yc3nIUtAgnTmR6WGy6u4KaUx/q8UT38oD/keeS5d6fplkasBnxgDJSN
f3hhcSrf2zSNh9R47YO/Ev1mVNmrdYWKCezVsD461j/vEJwZ6lC0L3EkM5zGWhd+8/qiLYDLtDrj
clidr1h9FoqCy3ejeH07ys9FS3eRFtZrapX1ahYTqyFWP4IFi5+B9sCl/DcAjj4qvVVHSGTDIdQ4
xdDykI2lTiY/k567I89xmmYYhVuqdifABwZkNd8Ou7jkmLUde5xsIY5LxwZVkBa+HLVit4gRNOo2
IJAG+/NShCAJy1PJsEPkZqQSgVSWYIfMWErXXHcBWe1cM2kIKj9240jOvmahzji9mf8N8FbbHy19
yaQpoLWHCKnLX+t68dSlSBxGc0RjQW4ilStChuwnrSi1fHEBWKUjcj/btSAJTuPta7+xutuu2xRJ
cKQnbnYAqvKPNa5EYplsLtFWBoCLZs8FFpdmxZJkNVFwJzvnuEG1FJZSw94PN2h2mJu7frT9ee6m
6h4Gn3/RYiAeTDQVAmj/Qjuz2b84CsAOjEvMm/8M2xcSirsIN00CaYJLgCa+ofmbAUjM88neP1X0
o9EsQdEKTUYGznCQc0yGmML/M2J03qFlF6IAxeqaz+LTH6a4Ra6r5to756YQ64NleQjXDON9K34/
KnkSPw0LPYRF6x5wMsuKgdCilzxX+OzNn3pFwCVj3JNOcm9tEPg4zBGOitmAYPQVSF76w8f2NVyG
wkpqWOtPtyelFFlBSEW9MA1uU/YHCeuaZEU0/wKfRRC35t2Jb0mchBdI+Eo+aUZhFC2VugEUi5TB
kgjYWGa22NnB/ynnQJXTHrDuLGv9kMdrQbxXRsVeOEslwP5sehOnrToYJGfUagcqxL+eiuVTCEgg
cd7THDuCw5iZYVQoN5l4PgwFEEmmFwV1aVfW3W4vtj1tNvq0ZOyxeNdpYW1i3LYDo4XOYhAAxTY/
ms3fzjTnKr9Fe8gJwj+rEzSbK82jVghiynUt39+hNObOz+4FtVGGS1Knyv4JMJhtTtsggWi+kf67
BpwTKdndb7KnYdqdqgW2H4hTwDA8VtFrBGUVElsfKHHKI8THZdLOsXhxCQQGTHcJ3HLJijXbRQoh
KqCSHLOD0MlFeFUnvv0EZSXOv0UcSNIGIEN7H02bej50dGzOqYUkW9HB39BziHzDRYPlxF96U2L4
XDPvDBaMTFRQjEPXheEdKPcvBqS0QmZYf0VVmuOwfK8jtOc90j6YHBYpTfHLN/X7/as6eIDNFUR1
70wlcumUL0b/URK0LKu+41HG9CJzsR4/vFYbyG/4CmnUg+sdOEf4LQxRJl0pDhhV7UtxmxiA5r3m
5QjP3yla+r4Jg9Ta1ru9vOqJhZlB/LwMmbDF3hBtSgkO2LY89PkV1QaEGKsGRK8dlpZ82SJeMp0s
/tInGQupKL04HHA2sTaBfmrP749zOn8A/23DA6HS+2cOzzju29WcWitCgrkHND3MmEm60uFjuYHS
pQXD1GLiEVoC1cMWa5LsTbJ85NDGd72o6jQsGoMHBrMIT4aLAtHDOCR63vwitJBts05HSqC54ad5
IbynyHwit1bZhpfv77f56o4QnAcKz046CZ29JMtzV6+02QN6M+34eusVdPNqOhpldESkGQwnt7QJ
TtS40QkWY9CqarDQKXtRzIgPQqVXjvgJQ/2qJ4c4s5dq4AcSGAnb8HIB9o9GF+Ifbapw6LJOyn07
n+o8k/BApiLCcSATvnUJxAcF2IfHIOxbUijLDH1lQ0uEbUTLwzMwoH+EJG3/dqeABP/zo+N3/9ne
/R8htCxA44X5fjvd0JEr3kgTRc6UglSVBeC/Zrcn7UTIOjrF1H1Xe8dcwmkLO8bLqJ+Q3YDzqysW
387ekaZPPRZrU3/ta8IuAVpnPkPTzDVKH9oVdK0VN5Sj+PHwZG3IlH1pb5vt1qV8IMnuehPIZ0Iw
7Zf5UaBcYJ06Oh8ot7rKyFuB5GyjZum2LWLh4oSGBcimP6apjd577TLP+V6S1YVq+kyRGO+9mOBm
9wiovBMYy8gjm0/w/sH6MnysBfSx3Sozu9Kj75HQtPXEp5cjdew2TCw3RLPfMGLZasINvVDtBRKz
agOnlr7i1tqnRYtFxMDPOkrP18o2iWZY+vp8R+ru9/yaIFgcgWXv9+aJga6R0KXNBqDMVUnNXeqM
LDFJdp8kFETos743Q8iATVkgSehkwd+Ho10GfhRNQW4Db5k1+PMQAhM9mNhYM8ez+KdxKBSijLQk
f7RoSFhc4LIY3q7boxYZ+uN44n9SdzP/vH3U9ite2IwkdLQ+jevADeAW7UhzZMbI5xK89KjYGITH
erbvExJre4jTH3H5tlHeM/kuk2zXEgGUvvYP/RylLMPALs381UexKnMChKUKJj02juIpmoF3y7du
ZTVMU2DjnSfqXpMRcqMdhMXqlk3UHHqzsgiyg8MHJb7RmNxcwTalT74Sok76DYMnyPEXnJfRbrKO
5/SdirEmO1yG05MjpsO/7ueKgucP4bydDbx+QQb9I7kT9ainbe130oK63n6D1jSENhVD5UUhCUeT
9B9XxtrDSDdsLlRz4LDm4IRxyGjKk/+Zk7coK0V4Wc7aiul5RZz4ok1WlSC/erjNUg/QeLnrdHaD
aJ4Gob7HU4d/9tz2PWOQ7jHXSxIYdvF7xbv0yLc0cTSf5cY982KoRbHEY/mVUHGYZoiKYXzHCHlJ
5o5qR+ycaQNvmTLildXTqb/3wqraV2PWYCzeq8tgbE+oWx7+ZUhfyKETkUjiaXohRks+bm5c7Chz
q26ZGz4GxYUBhtAorPOXtfchBFZN6Ze4ptNxAjosvbpdLyqvHUi0jpr3Z71bbkjt97s30sbsPFsn
NFq8n+tWttQhSUE0xskKVKliG/w6QuCy4G9eZw1KHG8vLsnfsOPhwxVisbwyIskCKLHo7crznwIU
d5+7z5B3e6DOA3J1jaM1trrvUl4ZgiuCTnsuTttE2Z9G3GDCRSyJmdIiPTs7ICCQ/JR/4Ltbnkxd
dJbHhQrHFsnm8kWj+2EAAc9D/bSefkce3/CRM7C52ZSTOsPccokbk2H15Raad76k8GVMFmAIwC9s
PMJ6Z9CVtgveeQCJ6jvk4oot8+XNlczGiarM+nhtaf8yXQm4nrXqjP+7GXmNisX98hY+EJCShf+S
H+iqX2Ngmd9r9wou7aENz0QTeLMcxh6a51CTSgQeqM97iSC/L0xMD71FwmeWF2Ta1HrZC7CEF64+
67qhMQtopmFBLhDuV8ti8qZVLEck88B6VW1In9fV5xms8VCCVaUh3T4/56VJDc2PU92xTGMWkI97
Gb68fIferztqfmL2ibBd0T/0mSmc6TWYdqS5u1Rr1b5bljtDcxg0wr7JNS4IQu+kUBRu5uOQDPTw
l2CUG5y9sSfDtFE7Tr8RatqpaQkzvVBGeoPw2ar5t5n4gCTNrpaA10jwKVJ88FudMCtXev+DJABf
wnLrj+51XDiLQVRCJzQ2+eQrQfMONwq/cotEfcFXBx/+KOF6rbS7Pgk187pNXeR0aBkJhjnnZfN+
/+5ToUoBWMIyUWSrsoUo9qEULbzeHjcbDabIEVGpw7XJkXKrNzjBKEZvXC+ukQh8v75+gkBFwJI7
d+utrMh+e/St19B3Pxo/17hVngFUEdnCiZLOPJFeC/ZKI9Nt4U7lExsX/fHIljNHim2n89GbUfch
V8nKA5vDvRjyQOlhOf/gLjdv+JuEthNwNRjpKZ8G8GoAZ2qBZZgmzYVeS2KbOvEePMO5KXQlO1st
sGpqW/linDqvp0bgfAoz/UO0pLld7gaoNbUEQbGn9Id7L70j9/AF1T5fe6J4iIbvD2Hdb0sJOq7U
4/6EUJOijOEiI7DFtEamR7EGJPTWItvBHOwFSUfm7ptyMjbwprS+N9pJlYtEzuYjgfNO5baNjpIS
Hw5F3AHmbFBrX5xHdvseJ/L1aS/H9c1jLPNNKRMBYPNOVFOoB+rDeF7g/IjKF8xUFr9HtwlLBcd4
RnGVH2AnqtTCnSzchLkdn/tbumNylf5ERZFBhj9n58SST14pfg0RscSbCrSmgtYnsNoFd05ppy89
6FcrW3YpmwzWL+WCCTAV/HI7wMvlLigJr73+rGa7pIr5/HhsY54JE4aPg2aIVR8j4nHo53uhqwho
BISk6Whj8FPjVzPUbdnO+w1l7wmtoELedmMemLky9L93VLD2YP86aA2YFEYmnBIIl8pZMufT4nCt
W3+qnr8MmrOOFG5uTEQMEO+NRClO7AoDiz/bgwpb2HXy56+P4fp680ewgscTk8LgbkaRZ7H28EN0
uI+ZqVayFPYyK5sT1pcN/oRwqmYs6mQXqjJmOoPLwidIAD0dv+x2othGh+7T+c0KVn9B9gxIjj0v
a+T4xDDrsBgo6lIZjP9BGgb6s0msVuYU/SkIcNUn5XBvS6McYHGXo638rPim5cdAlJbdnAt+gbZX
g03PkPxAwl2YpQHbm3f5/HcrBngeGIDi+wOy0PMDYBCQEr05pCE6D1FpRE0KhzBAgibIbmPLa571
sXkxOdAU/0j1/+KQ0dH+0xn3CH2x11/8l1JBorBd2es/OLzKoj7MWYWM8KSXFPWskHpca6xpK/zn
Vkl4RJfUf9OuDmmBvV9ICacvdWUGkM+My3525tC/3RqDhkrTfsGxKG/BFCZ3UE7DYxx+OHE26PW+
FEzn79ohWPmtWZF0cbbOnvwezVAgPkByQ442KZ1/SMGBvk+US7WCmmIZrIcDjok8vLlNwosl5Sbg
i55hUwnLwSOolrtXCigLc6WR7o9jAHiq81yuOoG/eBEWJ3ApVv9MNhhiFNjAqaVYR5TWNxuejxv0
NiKUJNpapR3NX5GNlnkyy+qZ2L8rh08ZOuZ3OVBAFETGcLhZz474ln9TbeRsddrdiz4O0P9FRssA
ZGyk1ruIBlLcWq/F+wczcEW7lRw4nAJyWCCuHLYIY2uBOPeBhRUBo4tDkfpngNZsnkvMNv0COPTv
8KowHH3pln9YllPrSbVxZtn2Jmty528kau3+j2kEZ13X1cZBfCTe0gli4Md5AkawnsJPoNnsLAaW
LNfcU56eqpEMJzAP29egBxIeMehBWCGTka2meNvQO1JCTvj64WrtMXQ3I0HjsihspPqtb/gXvwhw
XXWQpDVSJI9n/gEXJlW4E0BqNUSMgzgCeOJkmyC57xoMFFjBe2DwWut/o6sfyk0mQ3aZvn2ze6ec
gZg/K75CUsdqBZxuZcPjccpEXoe/MbPp3MARXkh32oIiFDa6d5zhFqHVK/9cfnUm8X3df8iMlB5Y
s+XWnV85sC6PIyXJrqSxB+78Bn1T+lqvcOWXedm8KBFbUPh8tHZh9LEDy+CoJelw1La9f8JOeuBH
+8VtLMTZFpi9XOybn4dpol2MwvX9QLSqDeezX60pC6HKgM6i03W1t1Xrh2nECDPiDYOCYWQpFOng
LtUCewkK9Kit2mrr65JWkRvGA5tFbB121TtTJN2rP2rAZpcLZmmB655Z1B0SM0iZ2ns3ZxTyw8ZC
p+rLYSNr4p6+CxgeqocFeHpfAuD6ClF1L314JXHa86anZ7FOUl6TH1Wg4g3jf5WHMqz98bnB7Bgm
HN0LD9aDZ9+1FptCOyudopqQEJGUBsTjmASdINUodQmp6a1GrtHld52zhTopT88hS1nvp47/qwTE
+8kKeVq/zLpRoa8ZgcULeaQmgJpSDinMGkSVamlzlxHPXphutlHwXfPvo+sfoWCAzq5/LW+DZMDI
ii1+xcTPUnk7ValtRB1BoWAfcjhCxTHVIwApuV/ne6M3Fx9iCvh5UUHopT6mYgU1rmCLtDjBLy4P
n1Cm2AdzdJ0iNP/0CgzSCWAQQ/YS8Lk9/utxl/eV+O96R4/gpKb2ZkM56qTK2c8Pu1hBi8vJ89WJ
bvNIuacM5Y698pJ8lWCQC0i981egjNA12f3o7kYtyrtb+FsRU6/DAUx1Pi0UDDxqKs6HG7Bsqa8d
ugQ9JSS+9ke/GwiKeivnGGfDp8DuQYfERSi5pfHFOTGgXyDP7QU7IyahKll8U8jgEzga6x4fH5Tm
JjYxXwTVnG4VDtUW2+k65hzG6jDy+rLxeGyUfUOWVxFa2LioPcCQ3ZXFECSLUm1efV2n0CV1atD/
T5DxVd2RbzrhncxHqvntFD7jyWBqlS2+4CJ2fQDN3LqfO1rNoC4TflksSBWX6/LkKDqFfPcN5QNk
uQ6+d8rUwPaxYJ+iV0ZTh8WpTegOsyb7hBGXdONDLa6T0QhUh2uPSWk0OXYgNALVuzJOlbI1fcZ5
w7BZvxnivPDAsbJR0fSE4p/BNuch9ufCLkysdEY6PDZNyAVBEg9wTs4twNTTkyQMq0v5m9/k2y+3
+LpyFeEj7gmUZ7F08KuuuE8AoZZr96Bgk7WjJuAMExWKNCXEvzmGuYGKcxfYSWs9j8BoNXr9IE1c
icgErHXQyCQs+0M0vdWdTeuf9EflS/b1kJy4NpqDyHKkmuYqFUiqAcXikvd30xgvygPfk8NBDb0j
JsWYZ2oPKIswts9ab0K4x0X7OrR7pRJl3KbH8E2nIhqM9iG5q3md0X8jp6Q2sg7r9cZ/yEvVJay7
ne6shhaWsF+OhxhQGGRGmW+P/FDDPKPiGyLspJz72Z9cXP0PJcoZDX+coT1blKnU86g97/M+5ihD
V4gSvYuPTaaKkl6qzWvHiOyn/ZQ4cZDS4RaUOMoelHIIznTTh2pYJ95Icr5HGz1oXhSj/GrWZYcq
lwwYeHclG1ImhjZEmjXPqzJlhvOoedd7BtlPaEo/1uQiAjGenxp0dOlGIMj0K0iFPeZytsxZyrgh
xIT9eMd4AEEnP802BNwLn3TdkjfaJ9CJaOLYb26Xr4NW4H+8HXOYnf8iW76aFpcyK8IyMWutxXQw
PEGXCdFsmIDWzt7ycquCXBYH1GC/4E0DfD5bvdqxKlrZ10druAil5xc8bUugyLGTa7nWkbjeG1QV
RSnh0HmIJ6sHtOXGr4faJJLbAtbMNIMK5+UUdTqihJqoGtIVBIAv0PAdh6dmoKk0/puA3vDqoUEU
t60f0z/Gs4SrAxu4hpB+OGt8FlVCYG0HwRez4RzMhjN3thV5c6UQAEfxAgj7XP+olNwdkD93aM7T
q+itg/jxeRyHWB6bUxoABTe5XtFly9/nKzTgtllP7LXNM9fek8JVEXF/lCclmX2esKHcJW4FN4hT
JwCZx/aDkwphywKT21V13tMU0d7LxmNC+fkM1cGe84XPsASLMvke/ViVQl2cH/d3nmcOvtO/tlAr
Ed3nRLdw870hYpC6kO861nToxibqR3FQj1yUts2QSQH83ad+h37wZ303EUb3fPffTWUaY7/RyHqP
PZXwouUnVaZZn4XVzDGm2EHMLtTzpLiakl7OyD1+XvQx3kJdMLlQtDbL/B7goJGLRbt4/EJPZWCZ
l3+dobcKc5PvEeClmuSQTrghsve4XwrfWy5+a6bmngpl+bJseJkBF4WYXbyCdf6fRfXCxs//HYXC
J+shKGQhEOunNFf5HP++Sp+QhdqVbOBbCKeIkKdm4m8T5xpfIVLF2GeCZP3pbbX2kniAJpMyjqpX
t4UUlWhUa7Xs4jGSm/3bzUERW8Q3SvO3Ay8WGuawzpt87IA3n6PE3nqsA3FBy2ybYY/E63Fmnc+v
/HiP0To1AByb90PoNCYC8cms3goao22iTBoTiLSouI7UM75R6qJAwyoPzLvWB2TLZY0KIfAm2gmx
lk/5x4KucIit0QMVipq/2pP7pS+28s0HsxXGO0N10kxdxz7QN5xze00FvhddCMWe1chpr32ypZz4
EAMIrT0qhk/43q93HN7QwpYtZYMMPrzPIQCcp23m6v0vhdAOoJ5IMQraiHbWtoNy9FDp9F+srfIE
P+2sc6vi0y6zUFJE9nk0o0UZoHCkBZsBVXCfeizEqfxl/km3t1kj8Z6dIEAheqKF2Noc5w1Zj5gi
1Idq9LDGgqOAEyaAUVlXe4IOB3TIkdyiF/RD4K8YXRQg2uRE9dTZmUf8/QpLP3vBVQ1uGqghTEbo
Za4v5/Im5QKfcf/zXPn6oSCSefh9DeOgoMT7Bn0EeAZYqNpotAvSZ9xpP6NpFgVEC/taqgJrZBnB
v5zpwOh+CzQMz9a4UcmmOrQLQqIF+SSBDq3Nzb35Qhbr6vBidxI3wxWUFewSzbKtgHMjDMt8if48
qc16+oVjVVcYYGdbUV3by4jMWN3npVYLI9oFBB1xZPSezg8rUaPC/ds/oQUpUDhJIMvCvqTOml2H
BQ6SR2+/eO2wt5n0jv6f3Z7gyBVTdOox4wQZytIMl8uHi2zAzMTmYjBCUWnQUVPuhaeJaThYAmJ0
/H/peg88V0lxp4Gz7Ah1crrQK61AVlnu3GrWCYsst+LPezGoM8Zdt5aghDewsowuv4T1q1Gb19rk
Qr4ybytt7/Iw/pWQ82BWLGI9Lj8j3iiZ/tpmLmB0Ky+cBTzaCPgBAE1/un4ldm9roXusCk3UslHD
mPjHwdQDENQ3aGiiylB6PK3m0h3/b0pFLIkI0lnQRYhroUS8PgPI02F+EWDE3g1rYKomM0bRueBP
KRp42W/en4jIMV/ZSOaAd0qt4vwPixXA+yy6WweKrD9xkP7yIe2KUCNuVkhwHnoO5ecBY3yPS/FY
U1YQmTx1U/2/v4ZXENaISuh59xis9oBcUjdA2pxYeR/AKGUbagqicfYE4NrMGceNt61aB210aOP+
jJqP7hWkBPaRiBNUNz0LAs088AeCFHmU3Z6JILQ5Rtz7NWlV9oyIYuir5xGTiaJpA99HpCQ+slH4
cDuxyhBAraqXx32xnuOa5rnu8Q7AOcXksGcfsbIA4hNGTT4fbAv9qAdnS/vFY0IKf9MxRjzcmgTn
Jyu0/R4pGZKs4LHr2fMNn3tnIm389ANl3apLUPjMDgE2vunQb5XOazQXWfqf5WjXbYyjWB58mo37
kYfzJz08a9nRr6PYGnZ/dG5eFeqII10FVNc8QCForkwKtneNSkENl1s+syk3qwSsPOiBBS23NLGo
0oJ4xlGPRBz/glODc9oPK26v7jHXIxLULtwGigUpRYBUtwAJ+Hq1vz63nAFfFptkS8vpDmVsXINm
8q/SIyUHvDHZFrxaDZhadVZQPDUEUBh62l2EDYDZMq5BSOHj2j/TjhVMrWV9ecxeVRqvMDGn6uzs
ySCeaaMa9KqLGMjengu3tQiAHSRfY8fbrIlatY+xMj6WXcdoCxxyNc6kihSlB2yciU9yHY7QF24L
3MpNQLBSuCZGnvyg7oZ2G5dd/SDO9WwYFxn1qYeLf+U/p2C9YPHbrvO0Au6jwiGnUwT5mAgRKeNt
nocTssiViFCjMSs9UXyL3jmo+gc6+RWDitRLjqvOrFmm8Qn0O1r2DD51MXW2/+IvLCJqdUly9zjS
SMUiItHnOI+XWRcGAF9Dg8PdEYCQHPWGwX6Ff3mD4/4iwEhyye0OLc60EMaXVpS6yw0mABaNU/Xe
3bo+suwzCsCe7mOX98nRkfho8bzmf7SaDJOn6LJjmrWrAn1qrxfx5ilIG583wI7203YrN9cZAOlu
Q4b60+MT4T34AwvFHCeSswMloOsxiZ8ONtHRpLQ0OMumY9f08KXKfJuhrMxDSzC5t7p/VXODD8yS
FX/GbU1zL9SzKML6x/6ZCkFTtpd4YQtnhBUyQwq/vkQN5brhRyxGG4mX4ioz9Qdiz52H5Q51tr4/
QBZX+1/FxLBzHVGorLZI2bGQgr7s6wykyVmZEZ5nDBKeRPWI3HIplXmdXh6CkdwvkIu8aADmaTF/
AE1vyHqRLwK9Emi0L0J+BbxjaaLtpO1mpJWaLxYCqyOm2PsMkJ49nZZTBy7qYs3OLsUgkl742JUW
e7GtEbsLQB7iQNPbGYYr43oTYYZphfzEBVvGCAaOk6V7af+TGN9ny5CYBUUa6JNE+hySXIqoiYks
zgICcw8l9YTtItPuPLtIjiry4wuh1OYyzOGwAvZtbVbSvNc2HEZbNUWZY1E7P2mb1aKsAN/VPK/t
JNK/w39tnDSibhESrAHEzL/WE5y2LLdgNies1TAUGpOGLLJjUhzbt8w7NpjGKoGyLsmCzcuJTi+i
TclFTKTZZvxcmNQBPVJZm/PrM1SFOkCT5AqYRpII0ift11z6B4mCAvpNR6x54ICUiH7f//zpTPdL
8wyYZRLKO9XE0eDPKnPQgL8f6P9YKwc6AAbBu9JjcbrhgiROjiys3h/U1tRfexZSvKjHeYEwMiJw
7Wh/w5jDYCLYvZGGJhiFsj0XWlzFmlmFcAkwxDisg+S/ASckp6uo/bM1D9ICjoTXlcoqLX0LHfmS
fXvLn17TTBmD27elJ9ub3gcousac4LBNb61hDr37SUU/ZHllyrBlv0t7spOznT+Zyrid6iJJbN+k
quR0v2biD+JRFWbCm6Bj3ENgI6c361iY5U21blTiKUFtGJJQXU6Tsh8KdGWu6PQf0640Lt3Iaq+J
nMD8AhjRJ7KbVpkz1WFjraZ4H/KnrUxMCI1ufYQBvV8p9P+nKFeYJSnLo/BQbcx7cYXeiX4PFyz8
Mvxy1VE2gpcQ1aGG6NQacoALJudLj2hF/S2nFgIHmG/IV7cYRZUZCM0IWOJcHiCxgWQTBp9HZZ88
rOwMcFaLArVs0GO4v2d6Kbr9XZXwpd6C2n01zuLHuW6IslnmTsGNa4AvLpYYQwopHbs40QWJd8rC
U035LM929tGxaJdTlPwZ48hoyAHAoGolbGAuO307qZLjFnKA5dKsTbuf6p/wHK4T2wIgvdmC04MM
VNX2wtTsoowsO1h8DT7pLTlryZoYyQ671WwHptZHkN33SUbNU6LZJToij2YXhb/2Gwmm3JSA3Mus
uq5h3dpyn3qcCny5oJSIHR/EkY0L6DsC7v7FSLv+1LH9EC42BhU1d7HhravR5JvFN2OYcbtyb2+F
PtIEDmxRDXX2GNMdQnPZ5RU9dFENt3H/opGJVCvM9DbIDQVjZJOYCVpIAjBhkQQS+KAyllFX5Dlt
I5Dgm6CuLdafrzGO28/NOjK+Ra3AIhKR1v/UsXMrJikbTQ0y3Cqx95GBDgtu4KknbsWnAmDNQ/sf
IoIogeMJWvW3ruqfgTzKy/VkSBdTrczeWDFybAplhMgyj8hr70l/COz0rnykG+RgOBYjJGoe0wyt
ATTf7lu4EZUhTRl3EOfEC1m8xzeSfeE1rw/AXTqdBrH1fOBo4u9Djd8esxa/m57oioJvMTSVrJS/
9jkYsIcI0Nt5GY07WnXiVY6WkwtVQWllXNqJpxpwcFmuHUfo8SapDzTOgYmI2WEvMNigw+BsJJsI
44u+3rizNJGhqgMRsAFojF0Hw4yswrAuvwzjk24qHUo+leW+c1r1Rfsa63FMWIRwi4N4Y0BbGIkG
0Tl1bn8U9usMsCDfpmrRrNT+pTFzlxF7BM9ahSCon6uI5i8M1KgN+POALe6LqwCpY0PqFzWq0Qii
mgzfr8fHUCm0NhjYH71FY+2+6RESx89BjiJDSeXR+TaiJDZFX48zYT7cFlI+rOvaVlsvDYG399b0
rtBPgI0/aMssrdx6waARLX9PWZeZRBXpFqJgFqeBGU2yFYEYd6uuOLnC+/0IgbAonouJXbWDAf3L
b2EL0qXuJfJcpSRTT426NH6BV6U8yV3GHsbxtivGY+aDiiag6H3X79kY66tqDr9E7gO0JcDJNF3h
B+VtlqJGJi34+I6f+ZYUbo5KjvmcE/p3hqB94VslFfiIS4Xlf42+dYNYF4InQpo6I1igQiXiKEHl
jLu8Ie6dqOVMqZI7KV8/P/Y6fy9VrrGhh0cXT0XpCaKC11WechZm9+VowGpJbkkOGQ3hxvW4VKbU
jA/z5uX2V+fbvMMVYg3n2fe1FAOZ1aSadjVz5FFb0zDoJHZmtsP9JBKi4txy3Qg5kEBC30t1hS4A
uHvtyR1uuc2+NaHc7kiX8oPB99rY2uJZIv90yMdKRFKSCuk1z3jxl/yxU5Uick4U1yb24LzadYgO
2Ab0GNEb8YgCjr5U8INMYVkwhooQAoKH2jbEMJL1zzI0Z8bSPP0xcfTGgG6PCjhuLlWcv2XC1BDq
Dumf0MQefnvc6n8LOZKBT6L0IA7AVPecBhCauWZCunaRiTLDsbnwt0seQUJBTbKqutm4oE3hWff4
Hor3Pfk9fsCI86+P1IHBNsc963HlJIoTTslmn+TyOonx+Tl0LKzKBWgLlRnLwbdMKTa+jGqN4B2j
fuPFkGuoqErl6mpR8ufYXSqJ8Bv0Gb5KoSEOccBA2tm8wH71FouYsOQMsXQVIo4CQljDtJvi9XCQ
p9IEYO7ZlGbdzbmEaWHpsDNZx5HpSm12TCLJV79xU4iuuowsU2eRIY4kxcsN4ipAqvZVp+7SiFVv
+WtAVd1kxW62fgAZGNVzCL5FLrKAqNfH/9G5YAW940rqCtnem39/XdUXPt44IbtGm44I0iwjSjed
qheSm69MS6YOhOjQkDEMoXCPHklYPUX4LoQrMBk2C1Frg2tZ3C4eFEcbynCFZ5FmMrT0QGHsdHRG
v1x2Or2S45DA8dAm5U0mw7M6KzoqM5Pez25EWiPKtSH33/G1kbiG8EXroVeH8S1wBJ2dRGE93F/F
ar9W757C69b13H4krT8bkcHl3DOM5cxjHhBi+Xv/So0wliPp8PWU+rxrGg7cSxWV+8c+T0gdlTKy
kMD3BHXF6Z/ugB1yTyn643J0U4KSyg2syJBY1aifznUTul5mrBY4indD+UKE3IP6cUMLrDXao1q0
z7wuWggyq3j3G9KzAeYxOuebFY0PnqwHtVfMaOx14hTnvZi6d2tgkUb0jAv0sLIbgO1QyzGM3+NZ
9F2VDnqZ9it+UBrnQdBDSOGNguwoNZkJRLczCcBrRWVOfg+3XlnMVkE7d5q5Ip9tI2O3/YNO3WvL
ozZzaqH+NFDrXa+jGFcdo7eKCXgE8//m+6omEfqpUCG4RexxBwdY43cuLO9cCwlOwEsOS4vEffDE
FpIm53chUbQK7sjIjU87719Le6ApIg8r6BdDmHPRPJYb+nCNl6ieMF3EwOUYnBRA7Rwx7Rn4qXt0
zabhfCJj2xCsqlDsWGQsuzpdu6qr6adxTSFfBJfzR6WkzbO+5sTpv7D8jvQlkYFVM8lyFINNghRs
+qkULAlExVcshUCH7O4HeAzFuLJc7D44ONdVUWmZ0cY1LkqY1YuEwMBP1q7WDU3S250utsuPIW78
+JD+HI8nABgJ1htuodlPnl1XzHv0DbxvAbLpyqEJ1YVer9/0IYxNXFqSi9DnQuy+CwSTp/G+dHmI
BWtNqfrmyVvoYdltDQu5DWnrin0Gb2IeEA8xDOU8DdwqXulGYm4liI93/Qffmx/WevcWcU0/u+ql
7oU4VimJfzIIFW0db0kKEP/op338wrS5XBrbvKxdgqBYcBUS0p82pTtcr0wSf3HilafEtxLkcYR6
/tBJsyT72QpWJzKHrQi8nbEaLkWfOOvTfFpYDRTNPicGZOfNnJuPuZeUdw3h2zqVxNAHWHXYLQkc
roe4vnn94OYiUOUNnzYDRG/4Oy2GjH7l69MjCdzKOU0oOMrYkMzIUjUZ/ZKtuq8f8+1nTFYjJTlV
oGUyWgWoLhMrvgCE/H9lR+ORQgnvnIA66JeDHHHVf2Ptg33YPWzeiU7y/dbyHx/QTwKt4ANIoGg9
PLXZLr8BF4ohEv1Z7aANnAE1Ku/Evv9pFdVwQ80Wmp4Fj5ZWtuklIRRNGqU+PtX+FKKTaEFAX2RX
KEq/oJcZ07x+ASY9jT1CxkAOiP+hfOV+R25pUGF8tPRGHE+BAvgz+pc2/Bmn5HMhh1k5g1DDO2n3
MBWFy/s6C7I0cgU4X0ti5ing6QAZANgLEFQ07EOeSv7iU5hkpsRy5RXIj7+q3vDF+sDZe8lwBrPA
zpTxFaWFdZVq2lXIdsmM+liNA/+tERDcxa6oZNvIuvc9wL7TgUryuspFqduRheNXrWF/8vUkff6I
0Ss7/zv72Iv5a9hYcv6D1hcl/69TqUVIIi8guDAbXCsNfOLOxxlZeSP0mAxK42hlFEcFNRlbyzQ/
KZnW1jPdu3g+h0CltTj1pqzzw2lV0lKrRnTk9n6+8gDG5JQU1hb4Ea63KZea7nQkB+fGkEwlKVLM
LSzB9RHdu4WWzv3gDuaRJn29r4qJnI9jVzpFRyyvdJqHeAI9i+3mDhCpXzQ8z73+HCVy3XxDCPBj
lb9G/Jk3yLilU0nJhyIpSTVkdIVPz2V9bfdTW/RxZkyLPn0+P89QJmuFS2AZjbsyr9v6MJY+AXPN
WOy5+sjPiX5aLY7je8pkZ289upSdPdjvwmLYPbDtBiJsLlzvrJyOAV70twAhxPBbOLleCiuvPKqT
57gWUGzUfOv7AIZBGVLMAldHsvdc/j6NmL0FIfcrUC3O6jyoumyQhrQrmGnIks6BQLvzxPm446QV
SPzEeAx9av4rb4N22O1LwFw+jAZ8ko6UsHsz80djuAeJYPc6OEy1eW3yVR0B2/4dAC9AHz041fdW
P5S2Dz5z9ii4hgTyuE7NUuWdAVQRkAYs8kpDF/hfWKP3jtcMyzrAvQMn5UZe9T/rLQZgPsjCej/R
oT7G9Zkwh//dy2dCv29MxHcoysUS/lRgkKOQdOKUbIfPT0fQxf4JqY/3XpsKDX0hdqxINUT5dnTD
bbY+Y1aJOmI7TsYt7pJMkoqhb0tdZzpWlOAtOQK4wVL3YjjJpAWdenxt037oxGfyEbE9729VNwda
EXeDUuACAYNHKCtjvwwpQOqBzarfCesZVyM6OZUH5ijmiQT2Bxop9J40LN/ScrGvXLdwjL1oNk0O
STkM5qQlVw4ZBVSyKdTGy9f68r+QwwQDOmUNIVrWzfRlMMsPm7/+jFI1hO6TYcodCGqxSUGm4rgE
dCQ5nE0HnJhkHntoXLS3MKaN7LBDJX/aGzg1a+1Uh+/8nUT0k3e73BUO9dCQLh9wwGBIR2aHi4rQ
BhtEMxFShAzuS/grrmUIoTNTvPPTap0QR8efNrx+1o7D6JmPwPyMwUHlj52MycdhLyVXkvRHKere
ZBU2XuXknZkIl75SvRCZkj2htnV7Q2KaDL5qgmrlv6/9VP89rZ4Z0q6WJ7oDTJUKHCRkJr02FlgV
HlnNbMB0HU/w01aaIaEogRtS2PwQ0f8qTkyoqRTNZYaThiC4Qb4GaYsYMJJ2eIvaNVKETU8t1dr6
Q6Pg2mHgu0Rm/4p3aw2WobNlq5fmRi8idVZfnpYACBUQzMIDxIu+9kofkMY8/oLVf3KTWjWXWsz4
JlT3dy6Bb71c+lT6IGIF++eWAM5Yy+vLs0HUkEV38OeFvZmTa1e2PSzpDcyO2UZohN6x0p1YPJPM
RDJtGN7GdzktLqrj+rR6vVotDh2fTdIfKLiXzD0hx+8NNAvghl7x7srd8P4cAsDaIY7iyuvwaRJJ
cLXGhU8+Bf3HCxyvkM14ZNjnmv6I2c6GwG5T48Tg9DsbDUTJtw+Ha0d6d7KgUUM2erFVxPX2n/CE
PYGFYkbVcjNaw0ep/LZwJvyDvPwHdokUmlDLutT8RTMBYFWNVmCB5Li9P8PB0Ga/j8T/FcQV6vIF
TCjeq8Dy3ifMLrNFnjM9FIjX1mjsbkZKPrmPht/YCXtZE9fZSoP4xZH6wFFvEUxl6Vjz+Y5D7Q2o
lu6xIpL3WDHPIATASISqjBnXnfW+5N6gS81C85uu7HYM6S/4Stliqg1zwDtYucJdG5ebikHSwnyp
0W6dHqCJBFb4/K2yTG4wCMsjsZaqIUAhWfbBByAQTGHCP9YTV3mUYt3teFj9CfOXYtlj1D2Cu4TN
oL6NL1mYgzzCbQcxUB55dU3AendL+xeOHmqNAkObuloezyHETkmMPdcnh+teT+EFDEIsmptR5w/2
SOLhjK3X+0+glvbk1JeM5XZFXFNulCiI4twAxQCgPDNeQn/5gye00pjRG7YFMzD2tVnaTSRlpiLG
m3Xu+Z9hGnzaXg+u+oLkH+L4jtCKGE0S1erxxjH4R6qwrr5m6iUnrtefr5aT40b+gCH+T1Y4Caoa
e/pd/UBhHLvh+GzFPeQ/TooxFcN9oAjDfjSqQv14ZnBNTnQIWkpdi5UzrcKBjcXprEBKVmQD7zYf
9bKJuTTNtgeDpi+jyTCe8KeBsn2dWPRHlfxoMsU39H9AAAHh+2oVxZTWFEyUSDss5VE3CwIXp2c+
ilkx8rVQqjVhZhU7t2KPu/CM0gxF2WeGgSPTlMYiGVqNbXsEU+wZaZh35lgsFYam+T8csr1BrdGx
BewMjHTkrO4wmkrsya5qGvkolHq7rYsaK0j/G7uqufO2aYEnFky89u3qHObNUrJdmyy++OV9kLGw
EfCBoopb+RcIjqLRhac32hyrq+8/6cPq6Tm/Bsb9UGg1Ug8E3VPBoyoFS/zW79MikeTSZvSVA4d1
KLK4nC9YjuRQSWwpANkdbVcpHGbUE6lK+szJdk8zOEH8s2Oi6qfldF7/nip3TcrmS/LHVfrkxiyN
atpJXCMx0YWBhG492u30cphcYUHqLzCTReXcMdJmPC/Az4WVxNPN4wyeiWxB6sygF1CqRpHhU7Hk
MHmXGcIog+aTY0x6n+HCwq4JuZodzSbCqUr0AJWOqSQZiH2kG5FaPIArZ3Wuypee9zN5MauFVBMj
FXOo8r1GDuAr6YxCwDYzfuTU/W/FepGfGc8rDLdH1mxdJnYrmBGGfzXLCMPVDCS6Q/mG9UX51h0R
VRmLL4GDTYeFCJCbJWLT1lb/BgRRZneNDD4wmABDiD96iBUOKMkgMLSfBC017OeqY4kk1TlpY6pW
uAlllHx0GlpN6cD8WpR8qGLQcjAA0EJZboYPTi2kD9NU6dWPla963mnyNNEg+Ah3/ESHGKr0AxvP
BCCwHBhPLZKQNvZg1KBvjWswmHV8lvlHx+qevdCLnEcAIzqcrKuXwxNMQ+6xnR+rpNSSVx67Bt7q
0hXhHCFk9X/PSnOTwBnsknJgxPjEaktU7kDXrZAPV9OX4GkzhU4CXzedJc2TVCjFeFB+saKlbPGc
Tanig9Puq8710pjOQe/L/7iePiPDCIHyXFTcEDiTZDv7DeClBDByasFCH79cndUE95mPqF+kEXBj
HPYnx/oaDAS4pvEpnIZf3riiC43ZFkRMye9m+RO2J0mfb++FaX7F1yC3SeFvkE/uBXx36rOFxohh
V9xqoQIFjrsto82+YUBBjYsBAKmt8Kd0DukJONGk1cga1L0lFTZRcI7dpyQglh0KeFSeCLl5EUUe
TbDctaE5BdxXMJibDPuOWgjI613Bn8ue2WR8pqS34QyW1J+s4vp6Ak7wI6+W8pEPG5aOWGUZi1Lk
Xer3giVrx/YSi/GhHY2LkArpBICDOPrFFqmrAxFSY4Ax+357oj9Mu0zLWa2KOXDhA9Z+z4mDWHoP
T+i9N8zM4eGDOx4EGSGuUCT8W3hu1eNHsOK1kV/gDmK+A3bFoYplSbKoN3KC8R/wZzROjmIyf8Pz
VcntB746EcmmnJ6tkX+GF7FoK4TyhIevQ5nV5UXP3Nxrlx0wF/beUlp48Bfj+o3Jlphn7C8TAC0q
uNYrNFj7d1RjefMCUP0orWbTqg8tqG+bPEJOqL8ONAWAklISqrR5lo8HnvYhqG5815TXOZYwy0Df
I8qTojkHw3dxZUXeAzFNwl7z56V3K8VahSdkiUIBwUI8cLG3oBH/qlZznD3r7SnCgqV51hBRRJR1
fFJTZ9CV8A22z9RxVju6K6zILKyH0v/5H0GFYEKrXriFIpkC7IjJBSmW0YP2xaQSobFaWWs7xQde
ZOzLSZB5KrJ8Vl3YwU5vpDBM8zinbKk7MFNUW/CzvmC02A9y7TLOVEX2YpBq7pak3ohsjmmplCXF
LWjTbftW4ZNswRsZsbB67jWQJnW7Jku5AARHpbmvXBC5JIE2uGCez8KtRhtE9/X0O5HPwOWK9hCJ
ebm6XnciMAKGRymMuQSLd+syfjN5cxc2Hc4RSLYZtn6xxv6TeFY0jxqRl6fTIXZnkNyytIv0THcc
6fePQH4WEGOqo+sHD+dnWaOM6MXi0z9SRze7tA13cxeHTDWluorNVzEIq9731Gy0mVCh7XnJsPpW
zYD4TUYPs2Bpbja4YVYsSNlKIwdvTWF8xe+xnei0N5/ozZm8Ra4qv2iC+scC4KqsLeHteGcGswCA
w/WQ83M+3J2vaeRx7sghd+68qZdwgL2smJxYXBFmGivJycRb3aDa9H272X4adqHaZCykiGC0fcl2
GDV35AgfmZALoV5zsFzzEXFa3vYfpgS8R12dn1v5BPYsty12oKhHei5vUX9ZN+cTi78KwQc/jdYq
Dzx51GkMm1ZDDFgeiZhbdg25TuxBde74uSHaYILnYE9cZAWsQ+BntlqEji5mwGAibHZG+hu1TOYy
YccSljkjuU848CN4nUBbdHaRHYaB1iTLJXZUbXRoU5LrwN4auua7yhtQsu7r+s2ApWmidNJGB4g6
FdE9eQw1iF6K9YsY4nm09yR5nDc3GYTyDDsHuRaSA4uWR2YwRV6zRCMCAwaXyTkgn+LhDHpZFlxK
H8MTjHjfUGKiFnzQMQuSI5+2s58cX5uci1EdDAmMTMfRvseJExERnskwXI5TE11bPunG2R8tuTpf
JZrIJhWQ87cpuytT2A6fL/cCLYP0/dVF6kVAS5vlyZcdZjoaeY60F5bpbHX6BkBATwxnRj3zvgnV
hhfq0P77+8FS5SQn9S0AAMCuOYC08nISbnQOEz1OV7GLnJQUjGnh98ACTkWKkNNL5KoRdhf5Jnn1
NLNQCkWEjH4s8TJHB171SuMHpmyE00Usnh9fM+ouV4RvJzgm5pHZ4VLb58Wv4X5wjS9Tes3NSzaz
e4TPkE4Q0kPBeQHWW9ouYFYRcdXju3z4PB8ATx1c/JfRfZ0/GtvOuR7R3X0yAsl/ht2m59sO8BbK
FIRBaX91YlC3Kt4+N/qOrmBaQooe/tRwqibeWYq/p+y9yWoDMtpuU+OQuMEhEOWNJAcrSRRZUbJU
w2mHmEjbHlXLGlgUclqyhJhF6ct4xlNAbIf6CF50NLXy1HaBqxNQq7QScBZ14JZkpIYczp3zZRql
HAvwe0n2ciRPbYkz/TNgqpP0UiEiG2yE8eWUjTeawwiKIl0kDz9HpWzsXpK2uBlr+aRRV/q0qMBE
zj2/qEXR6PccxlHBLm/zopm+pLsH93kCD8Vj994kVVO8webhhxNAbpYWuTx7SaJCArGQL+EFM8DX
qk+smFavrWd2cM11fI4go7PPKZ5BbdtRG5Ujrf6aZua/sRhag/WA+O9zbVZKIRdxh03g00ROmi1h
wdx7JYVIE/6ACd46Kl/GjADpbvSxWuuQd0sllksw8XI7gyPS0/2p/uLp/BHpg7TKDOwY6obXqmZK
YL662c8Y9CGCsjzuBwz3VgM5GbuZM2Hrr5h4c5Tyz0p8EwMxuReOAUGsbpiiI+wzNQhOkkHWG+6b
JtJeLu1UYSHHi7HnegpN3HHqFLLudd2Ezbep1p3DQfTUIIQrizm5pZLdv3PlVp5MsIaYXQc6h44f
IlUWVLTISou9Amp5OHe+4sDpAYaLO9yG0u9Z4BrQbX+2EoOiLBQzW7l1P8/O1IoIz8PiWaG7o6p8
V+ke4cTv1Qnw3nIl+jjffRR3XgvVjZHdvTKYq22rscLxd6wEnmOiYzFhKKwLPgV7dAI+20QDhxID
gw2QRMn6tIFpf6apY2k5BS4u/0ju4OdBc5DkvEUiJgNVjaxwLp0+zxB7lJE4zJLfFwQvDfuOAW/L
jhJ8sBVkLVPO2nAEFl5wCewlbcgRLP7LeRPgdnx3kW9eQUwpTxGuNW220IilD3+wwzzqBnbkFn4Q
9imR7Pi9Yhr2TBIcKEQ7TluupYhBzIprBSLgUIFE+oXR/yg78TMlFgi/ONSGuZWDqdtf4tYZQ8HE
9CFEXkDWlw5KTDnoD9BiKeUQDTbrlRqoSAHHGUw12tUkhQ0X1qTaFBIfdL1L8jv6mcfxnht/sKOy
wz1i2sl3RgyBuU7ufTHCRMPB7eu5lI4+gqVsTeexKCPiL8u6h8ExnLtsacVp6r7ZRP7lQ1iotl2k
n2PJLw7SsqmxvnXdztEvLK/ubeppmVC+SsgvuastXJ7d3eT/AXIJ36fIggLP8yuHcy++QA10UBlw
MnOQaDp4QI74c58mJuYn+QSbm9gDQw0Td3gSVOS0PXlWRghVJybf2uyVPiUHt1EOtrHy+5+uH3E2
7gqJO7xIUYyIiLhQancc3COQR1s5X1+DFlIrlFKiwNUZnNpt6YmRWdOEwzlCzJyu5nkLekU1YhbZ
B0GNn6uVYHMi0jabs0N/GzT9bIAmYOhn8ZQ1X3+kyRWG9/hReM5G4poAP/PUOfezgGyzcbVy7Q41
eZQ6+4Ipyh3TGO/hA6HHFVu8WxONOJkAugiL6LMiL7XkkIKQ+A5BG4q9Cwqjtjmxx7Belde4hZCO
J0HH4bY3Yz8pLogYE/jFdVhlZ4o79vrrtAW+f6+oTYkg2C9zRbykMEiGl1yrcWbi1XfalcVAS6Hq
JGLTDUVEudTH/PnpqQdDfXT2Om4Joj28XTIGBi2GJbWn+OXzOZiC9nR2bWkjClWo4Gl3uv2+3pB2
pBEr6wyHDLCpapDeHCYEzTe/J3Hqc+KM7+GpXy3l+JmNNtomHiN2noJnNnvBKXdQ/tt2R5Qe2n2h
8Y4ZGe9pAUZ1x+DSrE5nuFQVIXzfTPdNiWy4WzpwYiY9dURf+E8GOLBn4ysAC3NfIjlm3Io4OCWI
uhLIH9Wb8ujRWEmepkxU8bqAYeBjYQRm+jJALujK/bOSKu8u5wwLoNEA5JeXeZ7sI5HhGnekgHMr
9clezq5N5uDFVDwBLcSdHHjp0D3QjTkgwD7COdOSjfA+zB/MSp6L21NJswyv0YW0nz2fMDpiclO2
Urhg35Uq694aZqHUM6d2zOFRFSB7J+29qIW4Ix6s/X9TeHLxLQTi+m6dqpbtiffW/vnZ8DrpV1pI
PR67JLE+GDM/qNljME2fLwAEs+LXORm0sv9qE/ulsXBAOba2z/LDcvuteXcUMeMoTVU+9b4NLFfv
FDALX1uo/j7/d/94SgFQnth2GswsreWShbBrxaz1uMcKhC/RWMvF6NbLAS55r6ldWnh+CsG4BwUn
iT5GDLgKVkI/M7WUy3GDUQ1fO4PaPv8xfddhwfOa5Q1TTZxAXApEjdXaIzeP0FiCjyqB97AI/Dvb
/Z7m1An8vZQO3lj7qsmOarHlKt84XjB6hxM7ylWj5tFs39RQWBWxf+3uAnEKyPS57f4jQtVXsmrE
5Re50cqEXzZ/Wy4tNyAaGF+fHVB6vlJui7d69c2expLqKxZ6t42I3VKFF5oRSIKb+Zs3AlvhScLz
TFjCBywtLUAqj+23fNkcwLwytL+hgVHLLZLoIABF/yiR0g3EnTwwfJpqCkVwPZJaMvgCsSr/AUPu
oYGJtTfwCiriz0bgx7M4QySW4PeSiFj3VIDi3vcxLFNByK226YZmoMMYspixpOz1KZ93DxqBrfp0
22H7nIBxJx32iwatwL/tadIQvh9PV7HS7E2ns2ARhv+dfCjBvzSGlysVvYjFQN/RY+uCOHIaMSUv
zjdlNXYW/oxbERnoPMaitZZ86YXkUYV4Mn4imDA2D9ZGDakRY9Lpn8f47OMR/hxuBHQojrh0nHgU
zyBxyjW23jEKMVzA0crA/K2SDx0kFgL14HhiSCl8kcvBUBmNGmZLCGAuJSs0ct2rvU8LtADYEqdq
15yeqCy/+oDW03R+pRmLvwmw+vGI7ySCXaq8dMlXxUONLYwFjQYfaSD7DkD+m/VZnk8Zwa9HinEu
8QQ+Qh8m7lEInkhUbW8igfEa2bCf/ijLOYiy9griBx+RRlEtCKcCHICi39HV12l3VwqJ4qSghUmK
ky+p/SSgYZ95qp8gzHE7C0ThoHbdrX65Gt7ttGHLejy3DhWT3FTEi2nomMaOlBtwuHG1KwzMys13
ca3OX9nOvxLdEUbj1a0NzBBnEL7TGxfiaVUCsPVKg2TVbZBYGG+Dn69wUSrBQVJ0q61TFcz+jtGJ
5l72AJk0PcTRqVrYmnRISEACliIW9n7qpJJh+5efKscYjQ1e4pdeBD6NsJtDWlVTVlcJmldZY7TE
929Ub0VR+YgS1eQ+5jdfQqrZKJ9pxS3lwH2s8LD6nq37hL/OpH8hkkKN40pOLjg9BOQf5nJz0Wvy
dk2O9fjc3tuqAwRrLjgOhyryjRaUkoa1M9s1N5TCT/r5q1MEumvAKWOflFhwT3HmD0s4rgDxQDFU
/xKyjFHqpzanfDI2xZ+ppPe9jvILEEw2MuamwaXc15UKScp12QN1M3NOzhq1I6VEmV816hsXWCph
cjZy9z5bSXAJOFHf3S5EnVEah7sQpHfDHlRGdTA/iPpscyBe4lDyvfNGbCYu3uOo3Et69+pKh8ot
1Eay3ANBsLLoxszfqoLEfMAXz1+KKu9WQC0Fwph8TLUAQixYMNeZ+xp4X7CJqVkESE6BHuBJLRHD
9SMsY6XHNwAFAqpEEwtFwjW+8r/KOGcJlFqEKMOLx3P7jGQmad8GIc9eyOxG0eg0T5DblQUD/iJ8
/JEG9OHhJncCBKuzXWQnHpcOer+E4Xjfs+/KOxQ/rc0NAddS82gBno2N8jEno7n0lzkYqLpU6aKf
GiIUoRFDjoTdBE15XJidGbw7YWbuTtkO7tChjq/jIh0ms2bSnvJzbhH3bmv8eUYFC+wZkE8SuRxJ
NcDBZhsrpnnSv91U1u62zrHtOOy7mD0GT8s0sZX3qnBasGMO1/bHSMupTw5O2RZ1u1jlsA/Q8t8s
PLasiYWAodhtDmYi4IrAG2guOWNfkqJJYVcgiGdwanka3kPm7B3hs7/brJklOmrBBmxsZaYk9I+q
UadYdXZAzu+6XYIdcTs9qwLa8sbbLMCTy7AHVHKxAQrKskje3vRk2fIFycsW0vy9wv/IKbKxjnhU
LvPY7TDAzcDv7WmX/J+p6omDceV/VVLpY3j/EZ8C8E+IBhsDpYfSbnVI9sRpPdlcLxb86CJj6sx3
yK7ZL4hftsm5rSNPzjnzqxO9Ko5FDRfYZHlhWeTA4dJq2Dh0kDMNumtsdPTargpXhwWriG6I7MxJ
dBGsnqHiNmmeMnmWZ4/eXNAPnztpt+wGI/FoeCD1FSMgEakiNCgAz8aGAF8r8y5mYOe0P6fPUJKP
PQiT6O/fxpMPutCqJB6BH7QwicgAw70ZiJFQc4rOWAV6VkgMcnRbnpnT1UMvmNCNeBdwRTFvtrgu
lcZi1AdTfe73VVGYT6aPgp57rJS3O328lWqoZIPTsqIqXiT5gNB0L4W24zqOZf7gi3H3Rlu4jSqD
Y6my8pxPLFYmuseP3foNmiw+Zgew0sL4fxN3Swz8LyDqX5ntGxG4y+t8lsfXF5PlbxO5DR8f1Zgn
ps6jmtOp5fO75aIS406HM9QroqUOPubWbtUglqa8Nk5YcI20rLd5G448Gm3U+bYzLWBF8ZMmc5ce
hOsDtZKIKruqcBagT1gyfde/sEBh6MsrtutPGTIpJ516K4H7i0rmA4V2xbr7VwDoXT79RrhlsQl0
H6gsipc6+/LP4NK6zKvaJ8ZjQjVl9sRFZ8XVooqN6JArCIvz735jZt4mJRu/SfDKp/5s3Pt4MSXB
bxNQuxC+zNDFUhDnuFlOVpZjcCl9UyCzmx2y00m7himMOe9MG1ff3dCBbPGVO2GhqIWOAOk+er9v
OYlV5/C6lRpNogyfOjf/RS9GTooHBeK3HTpKwxxxXQDl2VUK3AGlMxH426ShhN+0MPBn/6tSXgAs
HAxliVHAt+BNkwrxUXsknmcH5NPaTmaAgYfGYeyDmpp6dlTD+h4pCPu9bU+zVpMdY71wM/skhdvj
jIR2aSm+YuSiw3SSt0VDA+uLyP5C4D7PpxrNttFZDJXA3h56+wiMSdDhVDtZHwaqb88DwoQ6YRjX
MP+gfetvBSzAp/nhfM8GFOuPyjBPY1upxU+eg45qPn1XKB1mRQczORLyfbVBCDOxwRC7oxQNXyjL
HHBI6LDR3VMIIq+Fr9SQz3tbR+Fmn5Fuq1125HVQerynTx6cd4kEKWzqebjvE3JSpiTRmDU4xJiD
EUmT/T+1rJMmcCRJY36rFHEkxfiXTakdU+8QfEIJwDWbZ9/Ex5ZEIRGUTTKwkQUVTNl8Dex+ZULi
G9GpThUcOHdZRurXfUaMlzjX2RgVdIGfD1LQEXK3C+ez/Stx+7oaGXrHuYQD3szEFwC8eOUQYJZy
+ZBobTCpbPHAK+XOS67jwi2PXVnhacoWF+9FLqGS0HYXKIa+QCvByiREa8ZgMrLOkqlaiheLC48k
LjAAtRILmRmD+iP1H9CjxoDs1AO+MDT/Xbu+NDRWPRU+jWGSxmXrBXpcUY8r6ttYrf2c9s+NQbVp
2/TgaCZE0p0gvpxeDCCeYLxt2GN75u8IhiwtNi6JJZNqGqipnsWR+rURpEmG8KZb3lWkS9ZjeN6S
gSqHTWS1eENAi1Xs//GpMfl1Uq2q6qUJELLvdEUiflOO20+jv2MtkJz/9nUzdmzDWnqyfhbePQP0
BUytSx2wBl8V2n/L0P3dfzdpSuqon+r0hj5bNusQ7OSkSeJIoMS2JoGaGyx65j35id9hFF8v9HM/
UxoruNfeowd6Z0fPWzpvICp67b+H+VwsV6TK4FJRhm9ksyfjb99o53F7kN8iABY205XIBgWFqdYC
LHQFw5amvCs884LOznSLLAziR48G9bHn/1wufD3ci2HxVvglSMDg4TTpfb7IL+cefUlcUy2W9cfL
jldh4wATYXmZDVfQ0xVtaZgzQbOI2lKwEufxvlX65OOscABnjZe5TJWwDUUdxgkhwmOxA4SMY+j/
SWzoBaZbbVuHbFmJjLGRnPpZJ70JYzbk99OfxlVwoNm1Tn9EMvFHcOH3dfHVMbSSPIngQ50FE6l6
Vn9+/FKsuYTm0qC8R66hf4Ao6mSiUw+PLtOewYhc/pfki/l/aDGO2vpdq5QLpyPdlvnul68fDtba
k+HeImRtpfV/swJeJOjJGc0eV/PK/T3k78dABc0tDmcWVtpSKg3UfMqLmUi3CcBIDJYkh297ESmJ
2/nRmkj6mp1ZuLdWGSR1Epkr9wPb+dnXmgNF636kvdyLMx3H7PhAb3gwyF8KB6hceddPqQC8WJYa
jIYO5MSszsEsIcN8We95V/plVc7f+gRlVOf3MCqeLtdQ05N8SM7H4ccvtSx22BSVceuGov7IDTO4
1INcCfhoSSbVsK7VcPR2O91ScyCDBZqFlu0OVFDVCTK1VcKhU4PhXVKdeC5CwXBUVunGL6Q0ixc2
vQsdYsi81pauF6lQQX48z9h1jS1vxPy6ElBqytiXUFpAPrH8/HCY6YzqiyfNTfJtSKUGvdt+eRi/
bIreFP+R8nYIsD86g0+f+gxchQFBXaHAb1ZbtquVD05ggasmeyhaR2da+z7c7dwnuyNzlpluILKj
qUleHyySiS7gg1mJIskvwpll1pViNhvZYElGWlckQBxocRXxBsn6gsSxYTqqqMkK71FomONQfUHW
8xNsXtCEn75xTsYDA6OKMmCaMaKiXLHMgo+qIfLvO/5wkz5a87CovZH9Rx4Rolyj7es1DHmt+YoB
0mwn25hdCmr0epKmMVGPqV+dIfHrCYYTfo+VU6IRDqj1Tgxm4hmjYvZ3CZsobMbiK9uvNk39yJZu
+Cf5Gmsc1XdmCMQ7U9evvplAmmVl23AKEWOX8ZzhE6YKDAimubHF1hMiwBEPRj1Mm6PBHdmf7nng
mP9F3DdW7LkHIfVxYxKFz28k5J64elu+FqdhjW7WLXmKZ2vXnsNCmmNCEQvads2ULstRoHsHnMQ5
vBecn7uDFVaJHd+fWg/nulnmLANTbeQ++N8H2tDDRvcE6KenZ09TX9eR2g/dQX21mcGnO6CBSjI8
W0zU6AKdHSBC+0B1k9J6WyV3Nn0VXJJwkcahcewDJDRh5My3XjYt3Ms82qRpCu4xz1qzEqDGaGTz
yeAHXjM5gFufVS6ymTQJHcGsH1x5DretyNoXvSlv3mJxXieYSqHadk0SitTO9DjEgtgOXEy0Ei1/
UCAa5i4/x6eOMMLlEMa5VOClNpk9r8aWWQlLOz5BhF0aYOmHyVjtnCrbOLNFMecRIAJnhdy532yt
/B+X7sMYgWz28nmwiXseaQciPyy9nM8qgfKT33ay340onKfKfPg55tnrKuF9ksdWAZ9UpNWyZoN9
Lb9qJQrZipQS+F7QRjClsfolrf+lvLbQeejFvHVtkY/AEe9T4Xt0jYhxAxzF6sDbEsdfTIDiT0P+
h00DnZbv67ffNcPL81f/RjxUAgQnmKU0K9pZ+HteK7Cu8L0fgClYLIbwhudY4M1Zbzn8+FJ3yGhs
yk0mwtnl5fDOc6l3fL/ci78a5mw85hCknSnn1cxHXCUQNAgy+M88SL0VGfoASqHhr30PneYPCF3j
0+sR6S1sRJka7juKlLdNOjGEQn9dZPS5/GpVlI26GBERwkCBzyjeqJyyPm5atYVd2D2ZOLbPXd/m
AomOoVmtfZSgDAzOeQF6PJRBPIiieXFIrJaTwA7gFCT0nSqBW17G9HnMOT6FDW7JxiKfS4Ocq9G+
EkPGudXDlQNAjGEgSQgDJ6l5Tv/GstAfoKkWoimEBusT7GqADim9uZb/h0z0vpSFNBuSeiE5oF8u
fT0b15PzwhNZDFdeDyAiOu7H6lgiHJYYk9Ls03484c/qq8WWvzlRvhNejd2+fTpvKT7HafuYN9Ln
La4Y8/H4oGPLd/FnytPT/mziqP5wy+KCtxI6Q3bLA58OyKiLJCS00Dnj/yYGB+VDNAyVBjVuxBJ0
NpIn1Oz6H8z/1a7Z1R9HOxTPiBhh8sKDLmt6SKWUTwVI5Si6Y5WIahq0syL46dktuoUvOZb7inmR
HOTL8GZkdnqBKy1tcbf+A4Fj6Web8GDzjyIfc5Z199bGlavfkgl8MEgukiqyAvTy9OmhEfKWlOUm
GCpVz5/AsRZMQaaKA4o9HbnqsTTaqROQ7oeTPFSm4qDcVQO3SvCnGDuPSpfXkOIFN5bLayvwlh64
ZymTaGOzFpn4nHEvVphbav5EYRHEeDpmXuOQ9JyJyJrUu1f+KVU2/5uiI0/733DsDp9FxRCa+eVZ
hd54155Tmc0dyCAqG3NklwwsQiJhUhZadlr2LseLiLJWC3W9QBTF2ndmfX6cRwTCCjvH6eeKupdC
SDTpbpiAMDoThT6JCtia9FbB3WSkBud/crtwkBMjt4kYPr6N9wbQd2iR19aNHNHqNj4nvMf0YLn7
+yfmEIP2lw8AGfHxDOMQxIWPBg1pxYo4JnFe7g7pu5AHMlncv65ZTFATUrwEsORPgtfjXXvxGEmh
gY6dFB0MU2ZIkobZPiltMP0029Sn022t5U7a2EnnmQWCOGfqF8FIIFs03d3Ihlp/PwNZB71yo5EX
RW1s05BIen6AOqvskiPMfQP4OvEPmHO9IrJ4YU64QHsnzun7PmTZoGvWF00L373txo0oNMVbaPzu
sTL2FHFju4M47BjoJEvYCbfPeNbmD2fETGxr4IXY08kGablIRrJTYF9FOb//UEN8Swdxq6uLBqSD
CD+LUuxEdry1Sy6/1PglCG7HFkSjOtHxeXqbvo34OebaXpgN+/djuavytQp1UNne+sd1DzOrbIfj
auudzIQsBzFy03Uo9hpEvpiw7/lZxMfDvUmZFzyiY6naQlhzYWmANVrodwj+S0ekfQpItFP0OKeO
GOr6NXdnwfSNW2A4hSmXWJzL0zp3DSbssO2S3UtHqnEpLJOhjPH+JwsOig562dYpGIO5OYUndoKq
ya99pvYyDx6uBxMGZH9kBxhT3fPACweQVOLb7bfSbJS2MlwFOsuHtY0j0q1/XyfQO43Y10rKeF1E
30s82rWx+2/Cls2wl0Jonc3jBnKtAVdBIhpmvJrzejqFSLt/EbHIzSd+QNUT70anNdpCVEtBde+L
0f1KZWzvsv+w9Prno1KgnA1fiAPjouiYtprwR+QkUi8KF2J9MZY3DV9UcCFaSxO5AcSS0DpL/qSH
hMMaJ8qE7km8Q1xzYXMRe1caPz8UXmRCgHNdPWKajTEd2FRG/vUv0EbPXa3EE/7YDh1k1qCaxxoN
PaQ5imhCUr4QCAnpoj85A8iw/p20ySFmHKAkEDX+5F6DfURi6/Cbr3fnCgSHG47nex9Sgd1s8fxe
ZZ75QIpxvN2Mi2o5KgYdoADqekRClR1L+ePKhPWldAvl4fQBM/jeyJVPpCydVafvui/HypQUX/8e
3FLnn0Qd8ddPw/n58+qyLn2+LG/nMqXwlz49lc3X1Y0munNiWIWuo7qTt8myAvoJW6A+gqe5gPxq
qkzJk0Q8znbCZIp0Vrn/vgux4YT0tb7TnJlAhN+WpuXRYYrtFXHP7AE6ZxYoRnCvcN6HUppajdYq
DAWZ20i943bzUs/Js8wyyTkKzGkZnjj0ACygGIiPlnyStMg7l8RQb4kASSfOpDkD97eEI/Xa94vj
zQfdYpFAq0TOtNhdOTQm0vZdcZGSbHGq8aKUWlYWkU53xm+JlJa7Sbt4/uX8wRrwZcIV8jsEBEEK
AupFYQ/WfqrqgsyCJixAVF1yzinxlr8V61zYA1YjbfPHjHxzbsDeha+XR1XFN0rppIfNavaLcpLO
RFzkrq8NZA/AiFlpWITcFzc76ORTUn3jePu4Nw2xHTpSO+uVaFhFcswILMYRwipVZG7nanjjvAb5
w/yll0fxxHB/kkzSdWgbhgUokwDvjyn8/hhFMa8+BEeKvhRJOOaK3o0SH5jjvHgTZQehFYyRvy64
nn7voYzlq+aFNNXqNREeHFcrmmoDQ5gqq1W8jeyrH6N2e1crc7Bsd/58pr+LDPXFVBvzu2Q2HwNz
62Ry/5NhS7gojZBeXSovhMHamN8sNFr7ezdyUdJ4GMZo2r0T45xM4HH8tqB8Yciydi0fsyzXLldJ
9JvlaZVaK+SPzFh7Nx001/R4ayUBpkWJjxp9SM8iR43XQ3i9Xd5twKOHVklOz1guFW5INER7hRxm
JV+5DoPdSJz/RttsgajyuLfp+D2k6ZIJhEugWHDyMVOg6wUJvV+DZCg7UBAv9MAVn0r9rgYsAk36
P9+K77P+qY7tusAh8nzbZb1BI7pVhVoMa+r5IOR3e5YjqX65MeyRak32LA++o59MpZlgIZFTiVBl
yesIqhOFidXNQM+YOeGaaYo1zQYL4S1znskLj9SCdDxkAL83Rsdwri4+31Vh+UYHgWs/uxym2CED
4eVakmGhPBng+QAC6q13OdIkEjf8xS3w7qIr0WJudbkOixvgOeURO80XpYoz2e1tLpzR0dyPExKg
h00pG7NmIeiHVdqWJDiLeDKIUarvyj7DuCRsiP6gYgZqzh6EWOWjFXs0iYXvmKgOzWZJG6fUf1p/
JDewG6KM7CZMQ0JKsLsPs558Lph1J39uri6gsk3SQ2u65EPFCnyJt6CHSX4t0NEbE32v+8mJOvpc
nJ5vTWZ1Kq3tuTdAZ6FTnojbu6a4/7fDX5EQtB1ZDwRqVUqCfTFiYPiP+iee9zAZbPO4WK9KSSFX
boLNDfoBdXGVW3+mrdJX3sG84h+mx8l40PQ9Lb9L7T1ospkUOYQu2iKgRlwYAm/yYk+JqDe+P0re
EOkATyB+HpI/Wci3GS05JOtZGUJdxGKnEeHmyAjAF7YWU/Hcc5rxj3BFO0L3MOudSfe0umnSf3ra
krabTu1PDkCyCHKBMSPM+/QcYJMbmCzL+cb/s+9zYP7sYneahpSKy7M6s36Hk4b/IKPany1kNm29
94coIFugaR8igIinnIap7xstbwP5Z/PWNoy0ayhuzjYxtCIXlXs4Kp1bWhvlhQ3NOSXUbDj+xlix
DMtbQh/OxCxlMASmxC6QPAD3Awu8kysYuJzxAVQVH34alDbEUkv7s+4DgZSFxt6pgw56x4kmKkPc
AxYeXSgyeZ50TvWnwI6JZj24h8ZklcwkoSG3WfjXVilA5r0x0DF3AJ6m55lrqEKToBb/t4Cj8evL
PeA+zrge5s6fNdVN1Iik+8mgzjBC5gpVc9PrScgP2OP8B22nEba36yXY994je1+fdxYM3pSVdB1P
Q1Y7USVe0D7X4zzu5IpONqvKPdHVfhMT/fgyT1acQCSJyx9kpwF36/tKZkx4fqmuTJ+VAX+PQg/N
w/is8c4ZwpGU4hUQ07P7paFK+bIkDU13PHmut8SRHYODQ0xzmrCVuLRBhHhwJgJm9nXdFunxHGC7
UluJaVlRwnQ4T5l4tURpS0YBJYE2zJ9oQadHe2CC2vjPTq3D+pgqY2HITDqxtDHiJIhpRxGe57WF
HdBp4DBpO+mNmow4T+3cDoXyVI2zDvstz5g/v7BeEYodSdXRiK3JlPYTwxsrtTyetU/CSz+M4QTX
nGJiryMcgFlW0FILopQ3VAujxAu4d9EkhI0fL++xRW9AVvXo2paBc7A1RRuMYcKsDCLbe5V4dQny
7FSm0cZB5tsHGHm7rD2KDyTjn+rXbX26hBYRgAwlzljDZFdX8qSrJ1MI/Fy1uHIrIbWZ0QzfsZLz
AkEYzXTLVbl6fjs7OmKuufBqAJMiLmsMaARK62qLXwBHuggzTESNKWpcZ5N/EWn3KEBdReHUeAtV
luEME9+WWC/LvumzW3i43M0qL1gs+OWcJIeEcWpkkVihRlXWoVrSDpOu6CsaaTi5/h/lxMIH8qKR
LVVneR8Yxg4qDlp/xZOOqcmknkML+Iq6YS8P4uaGixA79zS4l+fau00DYwKc7R1kRTvnzWXCuXDM
YsUoQePLjehQgFm2t4kXOuDRkQpKdNviLcnqmXzOoz4JeKamNQDB3AMKE8u2ni/wn5ekA5rMXz5y
n0SdANNwYGkN9eKZBJG860YmWvmreJi4rPuKW6RSam12WKOW9MLw34eNY0KamOIMhS/68Ke2DFru
R2pEvFRKFovUUZ3yUopq74tc3k6hPURhYXs/xgGrNXj4hzIedLOtPfsS1MIc04DaXnZjm2BtePnX
8IpBSvNeCZou2I4yKdnCS05hryna1qUZLgED1TayjzgIGD9sRt/FLcYmwARkR17XcQVJ/LMMkbYH
47xVQSeSWsaf7c4Cw0e4D+xD+YFYd7x0OQ8iGZQxQ4Y6/gTXiUFgv2al/vob/jBjPy9jfUVxB4Hm
GwjoF0/KxqAQCKez3D34gJGNCl/1k7FE4H1mfcOR9uk0nUou9ENhdQUBSN5JqyuU1TAah2Pc9mk+
fgXD6+D1y5zPp1PkqNgcRfowXoAbyOwJH9dAmGlONojDWtElT61QeAEthoP4UCI8R17vtdnwt0JX
J3OxSpaYMwW4SJP7RGQ9/ZTixqnx3EwYieF4U4lJfyhBMUEW+wt7M5gLJ0pspa1Z21q0FTe8ySnM
kS7gL6W6Q6AOe8fUAuZEbe9zKi+q02DNRKlJsHijISb4Cs6xrSaRFG3cRxiBZILy2idx1BeAyNUX
c1+RtDcaUOQ1rkkujZAwTOxjVZ3S1mDhoEEG3uZL07/6Mpayu8MPKISBjvVVVlV+HP5G0amIFJuK
EcQFm8KeRdAwCfivF4cgzbOKDfZP8H8SPXdf6+QRzqMppreM1RaZNvWqpOaEPOc6qgJ/xgAsR5WJ
/WW20Jt3btYJF3G6GVGdJMA+Ckw//UZp7jVWe569N7EGFo3Gf16eN/EPHoa+aXvcl3hlG+fRl1fx
WcqEquV08+W3lOa+vlc0EZyFYo/KZfpW8kp+n6VXqrPT6jV0VTWj46UmY+cnWFEE3DfaUxd49kBp
q6NB6kn+P632XpGXeveLWGc9NczneN6MPqo/btBTmHv9wfHLRrcei1RB2rNSiDB756C2219KKReR
uHY8KwzjslYGc6Qw3BNOMpP5i3908WLtwa9S1bRWS4ns/YyD+3wRNY1XZNa/YKSLe8ZGBC+TQOa1
TMRpyJbgJI3maGqbeRAzTbD6z3uAUMaDUcploK4Bbsgdof/7kcQgpQ2tAh8RzCvPX7CXPyYckBpa
1tY1mbiNWOoISkB146Yl4OpNX3ZP6N5G4LpaJcbkUpjrVLoS0QcCJrhW3k71xyD7zk/IksXlo9jL
ABHZo3DwJeW4oeGHURfyw4rA51VU0rFLELdJfD+B6nwMYSbdbh5ovRdDylAwqJa26053C7q02u5j
NPZM6s+lOXUpOFd/Gv5XqVwHNGxY0Opujnn0wXwP+8K2qnxSiep21Tr9FNu7ozGAjlUvxgjUHSm6
t24165WKf9/Fwpck7Zm8i0P0p1wixZfKaJbIKEdBWnY4Q9JcL1BF9he/5EfrmE6RuuX5NqzHeAOb
LREcbbHO772t6k87TXglKuGEmym9D4f3VEMGpW4xUtoKVoM/QIXYlt1F+ZjtX9ztIkmitidjRfYJ
o4e67lw6shtKzmUZD05BtjYYKp68sj4V47r9c3XZC0d6O6K32g5y7jvMZxO1pccrgW1o9LRQWD4x
nOAh72AAcvHQ0rB9+Kiz/Gel801+HEVaa9oQ4epIr5wwNzUHtZdFHOeD3xgkqY/UapSszh8gKNzg
8OgxsYecqMr+u7bmIbQuz324Fogptl6SAi2GHG8rXk/vN+6Evy6CvuqNOFHUFMqnOX45U2foaB7W
TUj3kO6os756laYfnLq4M9WdbIRdFT52BjnBmWpBCodsQhytXNuPEO6/lhwFAs2gSej9zmAP89u7
XoLcTzasVH278ZR2Z3XQXacWublFPbGett2zafNh1Eop+IdJjl9OEt6fjmVumPaMyXt02WJMRlZx
JKpn1kNwq3KorzFvueSRqWHwctnMVplWcdUA8f7Oe0s5SerS7lIzFddgHEsiyNBvZootE19w31f2
hUEHEUw2o+qmumKaxz73FnwE+agM/mnbNEwKEH3zlBCKBTz/DY+rIuKlBniZeZqlWdaW46Od1HPo
Pt2ETrNMGSjJLuhvnawuCjXtcNArhGLBpWSwZk/bak+5yx57GvNMjdGEmkxf7PFo0hfV39TWtZAL
0VQxmE8dDE653mPKMg0RHenvcZ7Ok/KVm6U4fwJzTTm+YW8rHKbNYpT23BMfn7AtYUZTk46/GB5J
RQdnGB1Emd2sBRGXVE1XC96+mM1fF5Pr31dcLt1+J1CX/WwyHEiPLyLe5INBR/lV0gFORyWBSU+7
A5CbMeJrw8Z9SnF4vLFyMNKUDmNIrOXh7UXhudt77OnJiEVEMx31YjwFf+KxA5h1d5dsKFsoE/EF
hIHdDKd/WvZ30rNGPxL5IDAzrcPytUUSScNbEc0lHmZ0g1oLnW7jmCyv0/EIlG1/IyPefBV1nWPy
QoTNEbsW044jLF3CLlvHt0V9qfhLO955p5YDiDP/OFQDP7ap0CksK+15OyZ4agmqAUk+ME9TONMW
d81DkSi2XIJl/JjVRbeYrs1voOM/Y2jArRTIO2FpVNvD76mkmrGeiexbtce6+8IdzrDPTORPU8Ck
5d31zLMEpZYOpd3/dnQLjyvMMiz9D2vibMbJ716+pvo3eSH230Cgws66+A4aN8TynxzSjcS8r7uQ
hdb5IE08+pM3j5AvB9cgFdGHP5lo5Pe3PWorllihPZaaCHf0VMXkHgSi6o49CR7+b0FHIgQh837T
mA5xe4JPpVP/zy2e5eXaqqrPMwN5Wck4vLMy6pAP9Z+yCg629s7hKysGklSDKOtZjLJ2Thc6Acx2
kVTPIiYpSHSMMklrmw4hXKRvlmGJj6NgDSCi7XdPXkrQsPqKm1nTQPuuyLcI037iwYaiNwX4wZ5+
28NCD0/U2zcVbzehBhGfOaWDrn25IhXaxy9kA4IHhE9DXvrVr9kCgLOWNIHe/hWrVoTDlBO4Inup
iEYL/uSxpnF+wDn9AU3zosu6BVy21ELLtEbxMCZG9K1BHvJtzuRMmB8xylObyNAvZfewP8rgj6UZ
HoSpKTnF/pehJ9mz0CFE3+VfonAMxkRsSOfe5YSrl0297d2wCjLy44Mup+VTbelB8y+jrGs8RV0e
+ryNpndUZyoZcN8bpuCF6VTyoCo10ixNIGYIbbP4Rg/RqmkMt/7ErYTWk284kJ3acuPjJOru1msJ
uf2aCH4tQA/TGuGmB0V0Ja/dXSQu3II2GnXV+wi+RN7HPrviuA0tC5XgopE55Vl7SID6TCzr43h4
MJcqTHIGDSKFowUWvEuCwMOS6QUIIm2PyhU8cjo+lDTxVrek+l4DHpYMRAN9Hs7dL1OEqbMvxHyZ
WBub2HOoNV4PNrmZj1j5J5Gpsq7xlg42dpY35iDTdxZt70/A9Vt9XiOciA5xn8PMTZoEx9RhtEGs
7wMk683AH/vVERIYgTAj8VWwIlxicxFOIVPsJmaGwjtCwnYrRIvj2dfQWGtHsCnNUY0VBFY/j6G0
D7swWuPwj3aMCtIfq8NbqH8bf/kNKGFHfq1rlLboCh7DSAfjLXem8f0mg7TbaoIaCnJVCS6ocKke
PNuHdFWre5akkd3FWQH5c+NGHMlkr1rkNwpGnW0YDdq4C0HC8GZ38yne0U6J21y+AxcTqTzSU2wT
jOYZYdm3I74o9cWYRltpqmXmC9L1DLlPdug9N+y33BaVbKQXeyha6xdRojwDQ7I3Q7yIzOom8psY
JSjPhNdRjoOJqovkxZVpNnox1j7d7c52hdhE9Bj5mPNA523j1ecnU/trtJDBLpndpNt4Q0NTLCBO
/j/jt8CDTrFNDf9qQphsVrLjorUupKk2ch37L1irBA6s3XuMxv/23Rj8rX46M6rbNnH0/ixPxbi2
FkM2wsUMQJAJVWFBNz3YfyJtQeWL0y4CmKXHgDpEYVlmBMVv0GA+2nMG69S3JGi8BiNtQlnqqDxh
Jb+P7I/NThyVZl+ka2Lrt2oaEmGBL+dc19EXGJGXca4DxxoftcDa9MB2zKWUFQ9BwWX7dCBgH4+C
kxszXhFvIxb23jMtZOZj66RZBv4QhcTr8s6vtgvu+aryk/6pE/NZEqlPfbDeQEpLYK4xtjfk6PU6
9qXS574FxwD9Dv/RQH6JVlKZXm3wecCu6iXeoX+fIdwonNlj9gs/oyDJSEetbqBeSv0JUNPv0D+c
CmVvAyic8sD6yqJOEJfy8Uj+HQWZLMFaGWTY8qkBc9jCfAI+7SGctisvbUEYS+8IWp5+ZekKj/cZ
5GCuWx+bv9ylHDm2LsM/NcRvD8mWJPQ6U3piEbday5MiUvGR1L5e7qWZXRS4KvbBh+SgwgKhnLw3
6h1/aBfB+K+vpQLhI60odYh0nu8jR6ByjlIPjHabJqG/UOcqs+k9sh1o2oftOnah5GLjyBUg8KMQ
OugA6QWe7IxuIXkhO5X+VepLAk7edkpoIscGGvsCo/7rtw7ZRCt0YZODR7gZd7OzH3OxHWIJ00nP
j3dtlkDGGX6QM1cdYqgaSbinZ7e5Y2fxS2s35GE/LELF7LcGKKtYS5s+btArshF1TAk3nl+XVBlX
UVX0VOMwEYiFGmAZz61zJfDS/y7fqRmnIjyzpTSU3xwp2+ZxaqJWjCX7vCiX6LRYRWlbhHk/LudV
3wLpxHdU6BawRCR7OtY/CxtEOGlbjuQeNKVZ67FgcDb6GxdyA1QMD6xxCZV3oxgENn2Dk/UvyYOS
rFT2EmdN7lKrCMhc+yvVwbfqt1KpfSSzJzTT9++C9uOfJSCRcfL7QbjuoKj4zzn11XKfus6iTQVE
lDd4mK0dNwNLSeZpwygPfUThw/4Py0VguhjHOlwzyhizaGLxwWjWfeKtmbuy5acDjzce35QFRkn/
R4vOR3VghJemVJvo/QD9xrAanKL0y3Q0HE758fUEeicPFlPy7CIQnyIilwAqpcDLgTToiB1X4SVV
qXrVBEuZA0lTU9RAAa1I1lRncXqUWQJpNiCac2QI4dgPkgy4PPSxmq2J8+7/2xah2veEXJKukdZ0
TnnPq08l1SEPyjXIJwHxAAhZq5mnqBYfWthVyg6qe1BY9Vutc2FzGHHIsawTuWUDBqBdwUObLWMo
yg9fWUmra8A638rNUEOFBuabrX9q/jzx7byPBbYZ1ACQHuvUjV+e565us8KqbSx2Z0BEQ2EqoubV
gtNBf2+qhjwBcVLYR2js5SLoREsGQOfbm+mQRO2jpQnm2lFpYENiKDKyvJckPH7OqyIR7fTGAUfY
xVhiTFjrWRP6yai4BkGFUhE30cCWl7ooL938RqPC9bY4VqfDh1q2BAGV63lJYLFMUnjQYM40wtt+
s33qyiYTzSLo3wmRmxZ/qf54mvnn875uGc94TO9SRgEtbjQKoZOSqQ5UPpBjBr7ET6BG13nRyRwh
tWwUh08eW1jSIL3e9JUebY8JpAb6EcukN6x0vrAu+1crFQ/bcuCd4/n2dYZLukS54mktruRiafrR
VnBtvQy1KFCYoS0IfplHQJoThWpjKlxgfwtgyDkt/Bfb7qZ9/S9AtTBpdHHLTQFac8At/j9z2fye
QM7zirerXGPjlKPel0fh+OfWRF9vbfuh7axldHdNlAO1+Xf4SoB2f+zHQrDPTec91CEwdrh70tY5
oAEVO7OFPxdFN3uUEAptELER6HCF286bO7WTAtXhHBWjsGmd+A9kMy4Brxyd4nAsJmUSdzsqHTMH
9GCsYWPwEn0OzaLmzU7m50TT9VYX3n+QaUWi0qARGMrAD/lGbCCZm2AhI9+e9AEoBjQnlcQ/iBIH
1PWviHPirMFh/0/VNoHMB9H3gpT5zl1muSFOfWjxlWE5G+xGG2Q7fXnXZL6f93319Q6q3fAsNLpy
X3YqUdYoyMtAyjyhYtjYanQZGdlavRVaovkXbJfqy2y+eGZw6LpDbZpJDb34SoQxsjP6InQpv1Xs
fZi2+A9RAS1ATVzQvU7+VepDL9UNPqTcNgeBDfk+659FinALZVcbRuBrj+pMbWljOBRFtE1uu+0p
ikF0WBTiqzavfteaemY5TUKU2WSEe7G12kkJgtFQSjc1K1GAV8uZpymvB4AT+R16rw8Ktzt5SGPX
ysJNV0P41JuVooeULL4/XILdEegD8QSe0ZOsWCTKAljo3TJCMnT7O8X7Zdis5Ts91xVLcFS/OK3M
p7XyKUuJo8PnMr5os5mDOdRH0SZKT0EAaFODLP8E1gJ7Xz/BD9maGm5UR+uv0yDshc7lSvKAbH2M
aDiZyXMHicpSJEr8Lz8PSyE0Z159bWt4K29t99LziOAojsAGJgOIHzmDyUo05x0SQeOIw5x0cvHP
7WMloLWPQpbamGToJoaab64AMhT1TFlO/LXVfTuhGWramm8X/5OhJwcXQeP5GWE+EX8gAy1/r4vl
niDcaKGad8Q/SXG469LHOhneaCbc/Unr6jndciRxNOLQPrdicOwLQeTcwOsYhECh8zGg+jbgFzvg
SeddyuNO76X6ASXTHFmj/LRTA5/NuH47H1ix6O7CQYUzymg10QRBruXkqp2ashUAmLgn9uyKumeK
CSV9bM2lubV9w5hanrzux0uAKwPcgHZwaCUeyrMWzjFWQNe8N/tkin3MrKs0yfw5jyoTyUvh58Yi
V/Kj/OfYWcxuEN/QqII1Kk9mbEPdtNdrHp2+TOfbe+NibtrjvdN2PLqWkbyfDsmFMjOIAI+qZ9Jb
apVczLBIFkS2VhdfJDYUzq+DzqrvjZpB9RVIEt72UMhTdIGxRGPTtaTvtfOL+6Kl3S9vCO5YNw5o
rn5evYy78OmtMZBbdn6X0CM9cXsRbC/LetieC4QGZHqqdI5PS0QfjDvY8Q5PZnLEPNeQDEc/hM8a
Frp6mY+FbhRA9CXSV+mpLv3Jdyof+8BIce7Omv+g8qcvArSkgj9IRPu5/RGxKyhiZu+i9i6x0IKc
JiffN1XqaywzU2qyGmkUhHeGv49vgdV+Kf18gD77Rb5XDSULewsWz5cFIS9APOWbqNrLDAhzV94M
wgvWApFitLmHP9JD+1G7hkSl4XHA6BiGjGRPlxe40XKvdTSBEDNN1slJAXezrcRY13TFmMrzmZJg
gX+OZB+Prh43EpvSpt+xX2zQv/0J7ZWkIiD14+DVcJTCkuEzgjFW+37DlzJijtSD5X8FzOeZOt0R
4IWD9oRhmDB9x41d5sT4PFReKR25EeC/YMAXlZKqVkEGkLn2JuE+rG4k/ewB1ykWOS1C34NeXe7O
sATRaNJkjhZSv8soLTlD3Krn6ZSM42uUk0hDeWZz2E5o90OIhQhiSuf7bNnMGH6OhC8Fw/IFJOtd
qaGL5p5zhsME0Ir0572JzKLdVa8Td4b5GQ0z/jYuZy0aVAwMSAGooM9m496iIpjXaOJRPtQaMbtK
5eM/md3BjYu2j6eU6aaPfkVXsnTX67LZl4UooGfDx1OdqWXNbRJt71oDtPM2+eGMCOEL9chtWkTo
+2xojjRF2PielRSf7NSPTOVPcJBaptoEFQfWBddWD4Mb+OvDuA==
`protect end_protected
